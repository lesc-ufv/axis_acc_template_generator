

module loopback #
(
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 12,
  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32,
  parameter C_M_AXI_ADDR_WIDTH = 64,
  parameter C_M_AXI_DATA_WIDTH = 256
)
(
  input ap_clk,
  input ap_rst_n,
  input s_axi_control_awvalid,
  output s_axi_control_awready,
  input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_awaddr,
  input s_axi_control_wvalid,
  output s_axi_control_wready,
  input [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_wdata,
  input [C_S_AXI_CONTROL_DATA_WIDTH/8-1:0] s_axi_control_wstrb,
  input s_axi_control_arvalid,
  output s_axi_control_arready,
  input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_araddr,
  output s_axi_control_rvalid,
  input s_axi_control_rready,
  output [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_rdata,
  output [2-1:0] s_axi_control_rresp,
  output s_axi_control_bvalid,
  input s_axi_control_bready,
  output [2-1:0] s_axi_control_bresp,
  output interrupt,
  output m00_axi_awvalid,
  input m00_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m00_axi_awaddr,
  output [8-1:0] m00_axi_awlen,
  output m00_axi_wvalid,
  input m00_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m00_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m00_axi_wstrb,
  output m00_axi_wlast,
  input m00_axi_bvalid,
  output m00_axi_bready,
  output m00_axi_arvalid,
  input m00_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m00_axi_araddr,
  output [8-1:0] m00_axi_arlen,
  input m00_axi_rvalid,
  output m00_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m00_axi_rdata,
  input m00_axi_rlast,
  output m01_axi_awvalid,
  input m01_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m01_axi_awaddr,
  output [8-1:0] m01_axi_awlen,
  output m01_axi_wvalid,
  input m01_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m01_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m01_axi_wstrb,
  output m01_axi_wlast,
  input m01_axi_bvalid,
  output m01_axi_bready,
  output m01_axi_arvalid,
  input m01_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m01_axi_araddr,
  output [8-1:0] m01_axi_arlen,
  input m01_axi_rvalid,
  output m01_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m01_axi_rdata,
  input m01_axi_rlast,
  output m02_axi_awvalid,
  input m02_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m02_axi_awaddr,
  output [8-1:0] m02_axi_awlen,
  output m02_axi_wvalid,
  input m02_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m02_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m02_axi_wstrb,
  output m02_axi_wlast,
  input m02_axi_bvalid,
  output m02_axi_bready,
  output m02_axi_arvalid,
  input m02_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m02_axi_araddr,
  output [8-1:0] m02_axi_arlen,
  input m02_axi_rvalid,
  output m02_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m02_axi_rdata,
  input m02_axi_rlast,
  output m03_axi_awvalid,
  input m03_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m03_axi_awaddr,
  output [8-1:0] m03_axi_awlen,
  output m03_axi_wvalid,
  input m03_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m03_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m03_axi_wstrb,
  output m03_axi_wlast,
  input m03_axi_bvalid,
  output m03_axi_bready,
  output m03_axi_arvalid,
  input m03_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m03_axi_araddr,
  output [8-1:0] m03_axi_arlen,
  input m03_axi_rvalid,
  output m03_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m03_axi_rdata,
  input m03_axi_rlast,
  output m04_axi_awvalid,
  input m04_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m04_axi_awaddr,
  output [8-1:0] m04_axi_awlen,
  output m04_axi_wvalid,
  input m04_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m04_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m04_axi_wstrb,
  output m04_axi_wlast,
  input m04_axi_bvalid,
  output m04_axi_bready,
  output m04_axi_arvalid,
  input m04_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m04_axi_araddr,
  output [8-1:0] m04_axi_arlen,
  input m04_axi_rvalid,
  output m04_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m04_axi_rdata,
  input m04_axi_rlast,
  output m05_axi_awvalid,
  input m05_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m05_axi_awaddr,
  output [8-1:0] m05_axi_awlen,
  output m05_axi_wvalid,
  input m05_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m05_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m05_axi_wstrb,
  output m05_axi_wlast,
  input m05_axi_bvalid,
  output m05_axi_bready,
  output m05_axi_arvalid,
  input m05_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m05_axi_araddr,
  output [8-1:0] m05_axi_arlen,
  input m05_axi_rvalid,
  output m05_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m05_axi_rdata,
  input m05_axi_rlast,
  output m06_axi_awvalid,
  input m06_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m06_axi_awaddr,
  output [8-1:0] m06_axi_awlen,
  output m06_axi_wvalid,
  input m06_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m06_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m06_axi_wstrb,
  output m06_axi_wlast,
  input m06_axi_bvalid,
  output m06_axi_bready,
  output m06_axi_arvalid,
  input m06_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m06_axi_araddr,
  output [8-1:0] m06_axi_arlen,
  input m06_axi_rvalid,
  output m06_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m06_axi_rdata,
  input m06_axi_rlast,
  output m07_axi_awvalid,
  input m07_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m07_axi_awaddr,
  output [8-1:0] m07_axi_awlen,
  output m07_axi_wvalid,
  input m07_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m07_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m07_axi_wstrb,
  output m07_axi_wlast,
  input m07_axi_bvalid,
  output m07_axi_bready,
  output m07_axi_arvalid,
  input m07_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m07_axi_araddr,
  output [8-1:0] m07_axi_arlen,
  input m07_axi_rvalid,
  output m07_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m07_axi_rdata,
  input m07_axi_rlast,
  output m08_axi_awvalid,
  input m08_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m08_axi_awaddr,
  output [8-1:0] m08_axi_awlen,
  output m08_axi_wvalid,
  input m08_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m08_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m08_axi_wstrb,
  output m08_axi_wlast,
  input m08_axi_bvalid,
  output m08_axi_bready,
  output m08_axi_arvalid,
  input m08_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m08_axi_araddr,
  output [8-1:0] m08_axi_arlen,
  input m08_axi_rvalid,
  output m08_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m08_axi_rdata,
  input m08_axi_rlast,
  output m09_axi_awvalid,
  input m09_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m09_axi_awaddr,
  output [8-1:0] m09_axi_awlen,
  output m09_axi_wvalid,
  input m09_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m09_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m09_axi_wstrb,
  output m09_axi_wlast,
  input m09_axi_bvalid,
  output m09_axi_bready,
  output m09_axi_arvalid,
  input m09_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m09_axi_araddr,
  output [8-1:0] m09_axi_arlen,
  input m09_axi_rvalid,
  output m09_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m09_axi_rdata,
  input m09_axi_rlast,
  output m10_axi_awvalid,
  input m10_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m10_axi_awaddr,
  output [8-1:0] m10_axi_awlen,
  output m10_axi_wvalid,
  input m10_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m10_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m10_axi_wstrb,
  output m10_axi_wlast,
  input m10_axi_bvalid,
  output m10_axi_bready,
  output m10_axi_arvalid,
  input m10_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m10_axi_araddr,
  output [8-1:0] m10_axi_arlen,
  input m10_axi_rvalid,
  output m10_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m10_axi_rdata,
  input m10_axi_rlast,
  output m11_axi_awvalid,
  input m11_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m11_axi_awaddr,
  output [8-1:0] m11_axi_awlen,
  output m11_axi_wvalid,
  input m11_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m11_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m11_axi_wstrb,
  output m11_axi_wlast,
  input m11_axi_bvalid,
  output m11_axi_bready,
  output m11_axi_arvalid,
  input m11_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m11_axi_araddr,
  output [8-1:0] m11_axi_arlen,
  input m11_axi_rvalid,
  output m11_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m11_axi_rdata,
  input m11_axi_rlast,
  output m12_axi_awvalid,
  input m12_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m12_axi_awaddr,
  output [8-1:0] m12_axi_awlen,
  output m12_axi_wvalid,
  input m12_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m12_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m12_axi_wstrb,
  output m12_axi_wlast,
  input m12_axi_bvalid,
  output m12_axi_bready,
  output m12_axi_arvalid,
  input m12_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m12_axi_araddr,
  output [8-1:0] m12_axi_arlen,
  input m12_axi_rvalid,
  output m12_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m12_axi_rdata,
  input m12_axi_rlast,
  output m13_axi_awvalid,
  input m13_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m13_axi_awaddr,
  output [8-1:0] m13_axi_awlen,
  output m13_axi_wvalid,
  input m13_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m13_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m13_axi_wstrb,
  output m13_axi_wlast,
  input m13_axi_bvalid,
  output m13_axi_bready,
  output m13_axi_arvalid,
  input m13_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m13_axi_araddr,
  output [8-1:0] m13_axi_arlen,
  input m13_axi_rvalid,
  output m13_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m13_axi_rdata,
  input m13_axi_rlast,
  output m14_axi_awvalid,
  input m14_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m14_axi_awaddr,
  output [8-1:0] m14_axi_awlen,
  output m14_axi_wvalid,
  input m14_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m14_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m14_axi_wstrb,
  output m14_axi_wlast,
  input m14_axi_bvalid,
  output m14_axi_bready,
  output m14_axi_arvalid,
  input m14_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m14_axi_araddr,
  output [8-1:0] m14_axi_arlen,
  input m14_axi_rvalid,
  output m14_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m14_axi_rdata,
  input m14_axi_rlast,
  output m15_axi_awvalid,
  input m15_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m15_axi_awaddr,
  output [8-1:0] m15_axi_awlen,
  output m15_axi_wvalid,
  input m15_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m15_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m15_axi_wstrb,
  output m15_axi_wlast,
  input m15_axi_bvalid,
  output m15_axi_bready,
  output m15_axi_arvalid,
  input m15_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m15_axi_araddr,
  output [8-1:0] m15_axi_arlen,
  input m15_axi_rvalid,
  output m15_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m15_axi_rdata,
  input m15_axi_rlast,
  output m16_axi_awvalid,
  input m16_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m16_axi_awaddr,
  output [8-1:0] m16_axi_awlen,
  output m16_axi_wvalid,
  input m16_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m16_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m16_axi_wstrb,
  output m16_axi_wlast,
  input m16_axi_bvalid,
  output m16_axi_bready,
  output m16_axi_arvalid,
  input m16_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m16_axi_araddr,
  output [8-1:0] m16_axi_arlen,
  input m16_axi_rvalid,
  output m16_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m16_axi_rdata,
  input m16_axi_rlast,
  output m17_axi_awvalid,
  input m17_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m17_axi_awaddr,
  output [8-1:0] m17_axi_awlen,
  output m17_axi_wvalid,
  input m17_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m17_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m17_axi_wstrb,
  output m17_axi_wlast,
  input m17_axi_bvalid,
  output m17_axi_bready,
  output m17_axi_arvalid,
  input m17_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m17_axi_araddr,
  output [8-1:0] m17_axi_arlen,
  input m17_axi_rvalid,
  output m17_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m17_axi_rdata,
  input m17_axi_rlast,
  output m18_axi_awvalid,
  input m18_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m18_axi_awaddr,
  output [8-1:0] m18_axi_awlen,
  output m18_axi_wvalid,
  input m18_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m18_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m18_axi_wstrb,
  output m18_axi_wlast,
  input m18_axi_bvalid,
  output m18_axi_bready,
  output m18_axi_arvalid,
  input m18_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m18_axi_araddr,
  output [8-1:0] m18_axi_arlen,
  input m18_axi_rvalid,
  output m18_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m18_axi_rdata,
  input m18_axi_rlast,
  output m19_axi_awvalid,
  input m19_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m19_axi_awaddr,
  output [8-1:0] m19_axi_awlen,
  output m19_axi_wvalid,
  input m19_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m19_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m19_axi_wstrb,
  output m19_axi_wlast,
  input m19_axi_bvalid,
  output m19_axi_bready,
  output m19_axi_arvalid,
  input m19_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m19_axi_araddr,
  output [8-1:0] m19_axi_arlen,
  input m19_axi_rvalid,
  output m19_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m19_axi_rdata,
  input m19_axi_rlast,
  output m20_axi_awvalid,
  input m20_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m20_axi_awaddr,
  output [8-1:0] m20_axi_awlen,
  output m20_axi_wvalid,
  input m20_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m20_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m20_axi_wstrb,
  output m20_axi_wlast,
  input m20_axi_bvalid,
  output m20_axi_bready,
  output m20_axi_arvalid,
  input m20_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m20_axi_araddr,
  output [8-1:0] m20_axi_arlen,
  input m20_axi_rvalid,
  output m20_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m20_axi_rdata,
  input m20_axi_rlast,
  output m21_axi_awvalid,
  input m21_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m21_axi_awaddr,
  output [8-1:0] m21_axi_awlen,
  output m21_axi_wvalid,
  input m21_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m21_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m21_axi_wstrb,
  output m21_axi_wlast,
  input m21_axi_bvalid,
  output m21_axi_bready,
  output m21_axi_arvalid,
  input m21_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m21_axi_araddr,
  output [8-1:0] m21_axi_arlen,
  input m21_axi_rvalid,
  output m21_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m21_axi_rdata,
  input m21_axi_rlast,
  output m22_axi_awvalid,
  input m22_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m22_axi_awaddr,
  output [8-1:0] m22_axi_awlen,
  output m22_axi_wvalid,
  input m22_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m22_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m22_axi_wstrb,
  output m22_axi_wlast,
  input m22_axi_bvalid,
  output m22_axi_bready,
  output m22_axi_arvalid,
  input m22_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m22_axi_araddr,
  output [8-1:0] m22_axi_arlen,
  input m22_axi_rvalid,
  output m22_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m22_axi_rdata,
  input m22_axi_rlast,
  output m23_axi_awvalid,
  input m23_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m23_axi_awaddr,
  output [8-1:0] m23_axi_awlen,
  output m23_axi_wvalid,
  input m23_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m23_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m23_axi_wstrb,
  output m23_axi_wlast,
  input m23_axi_bvalid,
  output m23_axi_bready,
  output m23_axi_arvalid,
  input m23_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m23_axi_araddr,
  output [8-1:0] m23_axi_arlen,
  input m23_axi_rvalid,
  output m23_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m23_axi_rdata,
  input m23_axi_rlast,
  output m24_axi_awvalid,
  input m24_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m24_axi_awaddr,
  output [8-1:0] m24_axi_awlen,
  output m24_axi_wvalid,
  input m24_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m24_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m24_axi_wstrb,
  output m24_axi_wlast,
  input m24_axi_bvalid,
  output m24_axi_bready,
  output m24_axi_arvalid,
  input m24_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m24_axi_araddr,
  output [8-1:0] m24_axi_arlen,
  input m24_axi_rvalid,
  output m24_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m24_axi_rdata,
  input m24_axi_rlast,
  output m25_axi_awvalid,
  input m25_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m25_axi_awaddr,
  output [8-1:0] m25_axi_awlen,
  output m25_axi_wvalid,
  input m25_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m25_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m25_axi_wstrb,
  output m25_axi_wlast,
  input m25_axi_bvalid,
  output m25_axi_bready,
  output m25_axi_arvalid,
  input m25_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m25_axi_araddr,
  output [8-1:0] m25_axi_arlen,
  input m25_axi_rvalid,
  output m25_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m25_axi_rdata,
  input m25_axi_rlast,
  output m26_axi_awvalid,
  input m26_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m26_axi_awaddr,
  output [8-1:0] m26_axi_awlen,
  output m26_axi_wvalid,
  input m26_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m26_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m26_axi_wstrb,
  output m26_axi_wlast,
  input m26_axi_bvalid,
  output m26_axi_bready,
  output m26_axi_arvalid,
  input m26_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m26_axi_araddr,
  output [8-1:0] m26_axi_arlen,
  input m26_axi_rvalid,
  output m26_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m26_axi_rdata,
  input m26_axi_rlast,
  output m27_axi_awvalid,
  input m27_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m27_axi_awaddr,
  output [8-1:0] m27_axi_awlen,
  output m27_axi_wvalid,
  input m27_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m27_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m27_axi_wstrb,
  output m27_axi_wlast,
  input m27_axi_bvalid,
  output m27_axi_bready,
  output m27_axi_arvalid,
  input m27_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m27_axi_araddr,
  output [8-1:0] m27_axi_arlen,
  input m27_axi_rvalid,
  output m27_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m27_axi_rdata,
  input m27_axi_rlast,
  output m28_axi_awvalid,
  input m28_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m28_axi_awaddr,
  output [8-1:0] m28_axi_awlen,
  output m28_axi_wvalid,
  input m28_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m28_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m28_axi_wstrb,
  output m28_axi_wlast,
  input m28_axi_bvalid,
  output m28_axi_bready,
  output m28_axi_arvalid,
  input m28_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m28_axi_araddr,
  output [8-1:0] m28_axi_arlen,
  input m28_axi_rvalid,
  output m28_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m28_axi_rdata,
  input m28_axi_rlast,
  output m29_axi_awvalid,
  input m29_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m29_axi_awaddr,
  output [8-1:0] m29_axi_awlen,
  output m29_axi_wvalid,
  input m29_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m29_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m29_axi_wstrb,
  output m29_axi_wlast,
  input m29_axi_bvalid,
  output m29_axi_bready,
  output m29_axi_arvalid,
  input m29_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m29_axi_araddr,
  output [8-1:0] m29_axi_arlen,
  input m29_axi_rvalid,
  output m29_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m29_axi_rdata,
  input m29_axi_rlast,
  output m30_axi_awvalid,
  input m30_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m30_axi_awaddr,
  output [8-1:0] m30_axi_awlen,
  output m30_axi_wvalid,
  input m30_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m30_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m30_axi_wstrb,
  output m30_axi_wlast,
  input m30_axi_bvalid,
  output m30_axi_bready,
  output m30_axi_arvalid,
  input m30_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m30_axi_araddr,
  output [8-1:0] m30_axi_arlen,
  input m30_axi_rvalid,
  output m30_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m30_axi_rdata,
  input m30_axi_rlast,
  output m31_axi_awvalid,
  input m31_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m31_axi_awaddr,
  output [8-1:0] m31_axi_awlen,
  output m31_axi_wvalid,
  input m31_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m31_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m31_axi_wstrb,
  output m31_axi_wlast,
  input m31_axi_bvalid,
  output m31_axi_bready,
  output m31_axi_arvalid,
  input m31_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m31_axi_araddr,
  output [8-1:0] m31_axi_arlen,
  input m31_axi_rvalid,
  output m31_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m31_axi_rdata,
  input m31_axi_rlast
);

  (* DONT_TOUCH = "yes" *)
  reg areset;
  wire ap_start;
  wire ap_idle;
  wire ap_done;
  wire ap_ready;
  wire [32-1:0] in_s0;
  wire [32-1:0] in_s1;
  wire [32-1:0] in_s2;
  wire [32-1:0] in_s3;
  wire [32-1:0] in_s4;
  wire [32-1:0] in_s5;
  wire [32-1:0] in_s6;
  wire [32-1:0] in_s7;
  wire [32-1:0] in_s8;
  wire [32-1:0] in_s9;
  wire [32-1:0] in_s10;
  wire [32-1:0] in_s11;
  wire [32-1:0] in_s12;
  wire [32-1:0] in_s13;
  wire [32-1:0] in_s14;
  wire [32-1:0] in_s15;
  wire [32-1:0] in_s16;
  wire [32-1:0] in_s17;
  wire [32-1:0] in_s18;
  wire [32-1:0] in_s19;
  wire [32-1:0] in_s20;
  wire [32-1:0] in_s21;
  wire [32-1:0] in_s22;
  wire [32-1:0] in_s23;
  wire [32-1:0] in_s24;
  wire [32-1:0] in_s25;
  wire [32-1:0] in_s26;
  wire [32-1:0] in_s27;
  wire [32-1:0] in_s28;
  wire [32-1:0] in_s29;
  wire [32-1:0] in_s30;
  wire [32-1:0] in_s31;
  wire [32-1:0] out_s0;
  wire [32-1:0] out_s1;
  wire [32-1:0] out_s2;
  wire [32-1:0] out_s3;
  wire [32-1:0] out_s4;
  wire [32-1:0] out_s5;
  wire [32-1:0] out_s6;
  wire [32-1:0] out_s7;
  wire [32-1:0] out_s8;
  wire [32-1:0] out_s9;
  wire [32-1:0] out_s10;
  wire [32-1:0] out_s11;
  wire [32-1:0] out_s12;
  wire [32-1:0] out_s13;
  wire [32-1:0] out_s14;
  wire [32-1:0] out_s15;
  wire [32-1:0] out_s16;
  wire [32-1:0] out_s17;
  wire [32-1:0] out_s18;
  wire [32-1:0] out_s19;
  wire [32-1:0] out_s20;
  wire [32-1:0] out_s21;
  wire [32-1:0] out_s22;
  wire [32-1:0] out_s23;
  wire [32-1:0] out_s24;
  wire [32-1:0] out_s25;
  wire [32-1:0] out_s26;
  wire [32-1:0] out_s27;
  wire [32-1:0] out_s28;
  wire [32-1:0] out_s29;
  wire [32-1:0] out_s30;
  wire [32-1:0] out_s31;
  wire [64-1:0] in0;
  wire [64-1:0] out0;
  wire [64-1:0] in1;
  wire [64-1:0] out1;
  wire [64-1:0] in2;
  wire [64-1:0] out2;
  wire [64-1:0] in3;
  wire [64-1:0] out3;
  wire [64-1:0] in4;
  wire [64-1:0] out4;
  wire [64-1:0] in5;
  wire [64-1:0] out5;
  wire [64-1:0] in6;
  wire [64-1:0] out6;
  wire [64-1:0] in7;
  wire [64-1:0] out7;
  wire [64-1:0] in8;
  wire [64-1:0] out8;
  wire [64-1:0] in9;
  wire [64-1:0] out9;
  wire [64-1:0] in10;
  wire [64-1:0] out10;
  wire [64-1:0] in11;
  wire [64-1:0] out11;
  wire [64-1:0] in12;
  wire [64-1:0] out12;
  wire [64-1:0] in13;
  wire [64-1:0] out13;
  wire [64-1:0] in14;
  wire [64-1:0] out14;
  wire [64-1:0] in15;
  wire [64-1:0] out15;
  wire [64-1:0] in16;
  wire [64-1:0] out16;
  wire [64-1:0] in17;
  wire [64-1:0] out17;
  wire [64-1:0] in18;
  wire [64-1:0] out18;
  wire [64-1:0] in19;
  wire [64-1:0] out19;
  wire [64-1:0] in20;
  wire [64-1:0] out20;
  wire [64-1:0] in21;
  wire [64-1:0] out21;
  wire [64-1:0] in22;
  wire [64-1:0] out22;
  wire [64-1:0] in23;
  wire [64-1:0] out23;
  wire [64-1:0] in24;
  wire [64-1:0] out24;
  wire [64-1:0] in25;
  wire [64-1:0] out25;
  wire [64-1:0] in26;
  wire [64-1:0] out26;
  wire [64-1:0] in27;
  wire [64-1:0] out27;
  wire [64-1:0] in28;
  wire [64-1:0] out28;
  wire [64-1:0] in29;
  wire [64-1:0] out29;
  wire [64-1:0] in30;
  wire [64-1:0] out30;
  wire [64-1:0] in31;
  wire [64-1:0] out31;

  always @(posedge ap_clk) begin
    areset <= ~ap_rst_n;
  end


  control_s_axi_32
  #(
    .C_S_AXI_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_S_AXI_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH)
  )
  control_s_axi_inst
  (
    .aclk(ap_clk),
    .areset(areset),
    .aclk_en(1'b1),
    .awvalid(s_axi_control_awvalid),
    .awready(s_axi_control_awready),
    .awaddr(s_axi_control_awaddr),
    .wvalid(s_axi_control_wvalid),
    .wready(s_axi_control_wready),
    .wdata(s_axi_control_wdata),
    .wstrb(s_axi_control_wstrb),
    .arvalid(s_axi_control_arvalid),
    .arready(s_axi_control_arready),
    .araddr(s_axi_control_araddr),
    .rvalid(s_axi_control_rvalid),
    .rready(s_axi_control_rready),
    .rdata(s_axi_control_rdata),
    .rresp(s_axi_control_rresp),
    .bvalid(s_axi_control_bvalid),
    .bready(s_axi_control_bready),
    .bresp(s_axi_control_bresp),
    .interrupt(interrupt),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_ready(ap_ready),
    .ap_idle(ap_idle),
    .in_s0(in_s0),
    .in_s1(in_s1),
    .in_s2(in_s2),
    .in_s3(in_s3),
    .in_s4(in_s4),
    .in_s5(in_s5),
    .in_s6(in_s6),
    .in_s7(in_s7),
    .in_s8(in_s8),
    .in_s9(in_s9),
    .in_s10(in_s10),
    .in_s11(in_s11),
    .in_s12(in_s12),
    .in_s13(in_s13),
    .in_s14(in_s14),
    .in_s15(in_s15),
    .in_s16(in_s16),
    .in_s17(in_s17),
    .in_s18(in_s18),
    .in_s19(in_s19),
    .in_s20(in_s20),
    .in_s21(in_s21),
    .in_s22(in_s22),
    .in_s23(in_s23),
    .in_s24(in_s24),
    .in_s25(in_s25),
    .in_s26(in_s26),
    .in_s27(in_s27),
    .in_s28(in_s28),
    .in_s29(in_s29),
    .in_s30(in_s30),
    .in_s31(in_s31),
    .out_s0(out_s0),
    .out_s1(out_s1),
    .out_s2(out_s2),
    .out_s3(out_s3),
    .out_s4(out_s4),
    .out_s5(out_s5),
    .out_s6(out_s6),
    .out_s7(out_s7),
    .out_s8(out_s8),
    .out_s9(out_s9),
    .out_s10(out_s10),
    .out_s11(out_s11),
    .out_s12(out_s12),
    .out_s13(out_s13),
    .out_s14(out_s14),
    .out_s15(out_s15),
    .out_s16(out_s16),
    .out_s17(out_s17),
    .out_s18(out_s18),
    .out_s19(out_s19),
    .out_s20(out_s20),
    .out_s21(out_s21),
    .out_s22(out_s22),
    .out_s23(out_s23),
    .out_s24(out_s24),
    .out_s25(out_s25),
    .out_s26(out_s26),
    .out_s27(out_s27),
    .out_s28(out_s28),
    .out_s29(out_s29),
    .out_s30(out_s30),
    .out_s31(out_s31),
    .in0(in0),
    .out0(out0),
    .in1(in1),
    .out1(out1),
    .in2(in2),
    .out2(out2),
    .in3(in3),
    .out3(out3),
    .in4(in4),
    .out4(out4),
    .in5(in5),
    .out5(out5),
    .in6(in6),
    .out6(out6),
    .in7(in7),
    .out7(out7),
    .in8(in8),
    .out8(out8),
    .in9(in9),
    .out9(out9),
    .in10(in10),
    .out10(out10),
    .in11(in11),
    .out11(out11),
    .in12(in12),
    .out12(out12),
    .in13(in13),
    .out13(out13),
    .in14(in14),
    .out14(out14),
    .in15(in15),
    .out15(out15),
    .in16(in16),
    .out16(out16),
    .in17(in17),
    .out17(out17),
    .in18(in18),
    .out18(out18),
    .in19(in19),
    .out19(out19),
    .in20(in20),
    .out20(out20),
    .in21(in21),
    .out21(out21),
    .in22(in22),
    .out22(out22),
    .in23(in23),
    .out23(out23),
    .in24(in24),
    .out24(out24),
    .in25(in25),
    .out25(out25),
    .in26(in26),
    .out26(out26),
    .in27(in27),
    .out27(out27),
    .in28(in28),
    .out28(out28),
    .in29(in29),
    .out29(out29),
    .in30(in30),
    .out30(out30),
    .in31(in31),
    .out31(out31)
  );


  app_top
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH)
  )
  app_inst
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .in_s0(in_s0),
    .in_s1(in_s1),
    .in_s2(in_s2),
    .in_s3(in_s3),
    .in_s4(in_s4),
    .in_s5(in_s5),
    .in_s6(in_s6),
    .in_s7(in_s7),
    .in_s8(in_s8),
    .in_s9(in_s9),
    .in_s10(in_s10),
    .in_s11(in_s11),
    .in_s12(in_s12),
    .in_s13(in_s13),
    .in_s14(in_s14),
    .in_s15(in_s15),
    .in_s16(in_s16),
    .in_s17(in_s17),
    .in_s18(in_s18),
    .in_s19(in_s19),
    .in_s20(in_s20),
    .in_s21(in_s21),
    .in_s22(in_s22),
    .in_s23(in_s23),
    .in_s24(in_s24),
    .in_s25(in_s25),
    .in_s26(in_s26),
    .in_s27(in_s27),
    .in_s28(in_s28),
    .in_s29(in_s29),
    .in_s30(in_s30),
    .in_s31(in_s31),
    .out_s0(out_s0),
    .out_s1(out_s1),
    .out_s2(out_s2),
    .out_s3(out_s3),
    .out_s4(out_s4),
    .out_s5(out_s5),
    .out_s6(out_s6),
    .out_s7(out_s7),
    .out_s8(out_s8),
    .out_s9(out_s9),
    .out_s10(out_s10),
    .out_s11(out_s11),
    .out_s12(out_s12),
    .out_s13(out_s13),
    .out_s14(out_s14),
    .out_s15(out_s15),
    .out_s16(out_s16),
    .out_s17(out_s17),
    .out_s18(out_s18),
    .out_s19(out_s19),
    .out_s20(out_s20),
    .out_s21(out_s21),
    .out_s22(out_s22),
    .out_s23(out_s23),
    .out_s24(out_s24),
    .out_s25(out_s25),
    .out_s26(out_s26),
    .out_s27(out_s27),
    .out_s28(out_s28),
    .out_s29(out_s29),
    .out_s30(out_s30),
    .out_s31(out_s31),
    .in0(in0),
    .out0(out0),
    .in1(in1),
    .out1(out1),
    .in2(in2),
    .out2(out2),
    .in3(in3),
    .out3(out3),
    .in4(in4),
    .out4(out4),
    .in5(in5),
    .out5(out5),
    .in6(in6),
    .out6(out6),
    .in7(in7),
    .out7(out7),
    .in8(in8),
    .out8(out8),
    .in9(in9),
    .out9(out9),
    .in10(in10),
    .out10(out10),
    .in11(in11),
    .out11(out11),
    .in12(in12),
    .out12(out12),
    .in13(in13),
    .out13(out13),
    .in14(in14),
    .out14(out14),
    .in15(in15),
    .out15(out15),
    .in16(in16),
    .out16(out16),
    .in17(in17),
    .out17(out17),
    .in18(in18),
    .out18(out18),
    .in19(in19),
    .out19(out19),
    .in20(in20),
    .out20(out20),
    .in21(in21),
    .out21(out21),
    .in22(in22),
    .out22(out22),
    .in23(in23),
    .out23(out23),
    .in24(in24),
    .out24(out24),
    .in25(in25),
    .out25(out25),
    .in26(in26),
    .out26(out26),
    .in27(in27),
    .out27(out27),
    .in28(in28),
    .out28(out28),
    .in29(in29),
    .out29(out29),
    .in30(in30),
    .out30(out30),
    .in31(in31),
    .out31(out31),
    .m00_axi_awvalid(m00_axi_awvalid),
    .m00_axi_awready(m00_axi_awready),
    .m00_axi_awaddr(m00_axi_awaddr),
    .m00_axi_awlen(m00_axi_awlen),
    .m00_axi_wvalid(m00_axi_wvalid),
    .m00_axi_wready(m00_axi_wready),
    .m00_axi_wdata(m00_axi_wdata),
    .m00_axi_wstrb(m00_axi_wstrb),
    .m00_axi_wlast(m00_axi_wlast),
    .m00_axi_bvalid(m00_axi_bvalid),
    .m00_axi_bready(m00_axi_bready),
    .m00_axi_arvalid(m00_axi_arvalid),
    .m00_axi_arready(m00_axi_arready),
    .m00_axi_araddr(m00_axi_araddr),
    .m00_axi_arlen(m00_axi_arlen),
    .m00_axi_rvalid(m00_axi_rvalid),
    .m00_axi_rready(m00_axi_rready),
    .m00_axi_rdata(m00_axi_rdata),
    .m00_axi_rlast(m00_axi_rlast),
    .m01_axi_awvalid(m01_axi_awvalid),
    .m01_axi_awready(m01_axi_awready),
    .m01_axi_awaddr(m01_axi_awaddr),
    .m01_axi_awlen(m01_axi_awlen),
    .m01_axi_wvalid(m01_axi_wvalid),
    .m01_axi_wready(m01_axi_wready),
    .m01_axi_wdata(m01_axi_wdata),
    .m01_axi_wstrb(m01_axi_wstrb),
    .m01_axi_wlast(m01_axi_wlast),
    .m01_axi_bvalid(m01_axi_bvalid),
    .m01_axi_bready(m01_axi_bready),
    .m01_axi_arvalid(m01_axi_arvalid),
    .m01_axi_arready(m01_axi_arready),
    .m01_axi_araddr(m01_axi_araddr),
    .m01_axi_arlen(m01_axi_arlen),
    .m01_axi_rvalid(m01_axi_rvalid),
    .m01_axi_rready(m01_axi_rready),
    .m01_axi_rdata(m01_axi_rdata),
    .m01_axi_rlast(m01_axi_rlast),
    .m02_axi_awvalid(m02_axi_awvalid),
    .m02_axi_awready(m02_axi_awready),
    .m02_axi_awaddr(m02_axi_awaddr),
    .m02_axi_awlen(m02_axi_awlen),
    .m02_axi_wvalid(m02_axi_wvalid),
    .m02_axi_wready(m02_axi_wready),
    .m02_axi_wdata(m02_axi_wdata),
    .m02_axi_wstrb(m02_axi_wstrb),
    .m02_axi_wlast(m02_axi_wlast),
    .m02_axi_bvalid(m02_axi_bvalid),
    .m02_axi_bready(m02_axi_bready),
    .m02_axi_arvalid(m02_axi_arvalid),
    .m02_axi_arready(m02_axi_arready),
    .m02_axi_araddr(m02_axi_araddr),
    .m02_axi_arlen(m02_axi_arlen),
    .m02_axi_rvalid(m02_axi_rvalid),
    .m02_axi_rready(m02_axi_rready),
    .m02_axi_rdata(m02_axi_rdata),
    .m02_axi_rlast(m02_axi_rlast),
    .m03_axi_awvalid(m03_axi_awvalid),
    .m03_axi_awready(m03_axi_awready),
    .m03_axi_awaddr(m03_axi_awaddr),
    .m03_axi_awlen(m03_axi_awlen),
    .m03_axi_wvalid(m03_axi_wvalid),
    .m03_axi_wready(m03_axi_wready),
    .m03_axi_wdata(m03_axi_wdata),
    .m03_axi_wstrb(m03_axi_wstrb),
    .m03_axi_wlast(m03_axi_wlast),
    .m03_axi_bvalid(m03_axi_bvalid),
    .m03_axi_bready(m03_axi_bready),
    .m03_axi_arvalid(m03_axi_arvalid),
    .m03_axi_arready(m03_axi_arready),
    .m03_axi_araddr(m03_axi_araddr),
    .m03_axi_arlen(m03_axi_arlen),
    .m03_axi_rvalid(m03_axi_rvalid),
    .m03_axi_rready(m03_axi_rready),
    .m03_axi_rdata(m03_axi_rdata),
    .m03_axi_rlast(m03_axi_rlast),
    .m04_axi_awvalid(m04_axi_awvalid),
    .m04_axi_awready(m04_axi_awready),
    .m04_axi_awaddr(m04_axi_awaddr),
    .m04_axi_awlen(m04_axi_awlen),
    .m04_axi_wvalid(m04_axi_wvalid),
    .m04_axi_wready(m04_axi_wready),
    .m04_axi_wdata(m04_axi_wdata),
    .m04_axi_wstrb(m04_axi_wstrb),
    .m04_axi_wlast(m04_axi_wlast),
    .m04_axi_bvalid(m04_axi_bvalid),
    .m04_axi_bready(m04_axi_bready),
    .m04_axi_arvalid(m04_axi_arvalid),
    .m04_axi_arready(m04_axi_arready),
    .m04_axi_araddr(m04_axi_araddr),
    .m04_axi_arlen(m04_axi_arlen),
    .m04_axi_rvalid(m04_axi_rvalid),
    .m04_axi_rready(m04_axi_rready),
    .m04_axi_rdata(m04_axi_rdata),
    .m04_axi_rlast(m04_axi_rlast),
    .m05_axi_awvalid(m05_axi_awvalid),
    .m05_axi_awready(m05_axi_awready),
    .m05_axi_awaddr(m05_axi_awaddr),
    .m05_axi_awlen(m05_axi_awlen),
    .m05_axi_wvalid(m05_axi_wvalid),
    .m05_axi_wready(m05_axi_wready),
    .m05_axi_wdata(m05_axi_wdata),
    .m05_axi_wstrb(m05_axi_wstrb),
    .m05_axi_wlast(m05_axi_wlast),
    .m05_axi_bvalid(m05_axi_bvalid),
    .m05_axi_bready(m05_axi_bready),
    .m05_axi_arvalid(m05_axi_arvalid),
    .m05_axi_arready(m05_axi_arready),
    .m05_axi_araddr(m05_axi_araddr),
    .m05_axi_arlen(m05_axi_arlen),
    .m05_axi_rvalid(m05_axi_rvalid),
    .m05_axi_rready(m05_axi_rready),
    .m05_axi_rdata(m05_axi_rdata),
    .m05_axi_rlast(m05_axi_rlast),
    .m06_axi_awvalid(m06_axi_awvalid),
    .m06_axi_awready(m06_axi_awready),
    .m06_axi_awaddr(m06_axi_awaddr),
    .m06_axi_awlen(m06_axi_awlen),
    .m06_axi_wvalid(m06_axi_wvalid),
    .m06_axi_wready(m06_axi_wready),
    .m06_axi_wdata(m06_axi_wdata),
    .m06_axi_wstrb(m06_axi_wstrb),
    .m06_axi_wlast(m06_axi_wlast),
    .m06_axi_bvalid(m06_axi_bvalid),
    .m06_axi_bready(m06_axi_bready),
    .m06_axi_arvalid(m06_axi_arvalid),
    .m06_axi_arready(m06_axi_arready),
    .m06_axi_araddr(m06_axi_araddr),
    .m06_axi_arlen(m06_axi_arlen),
    .m06_axi_rvalid(m06_axi_rvalid),
    .m06_axi_rready(m06_axi_rready),
    .m06_axi_rdata(m06_axi_rdata),
    .m06_axi_rlast(m06_axi_rlast),
    .m07_axi_awvalid(m07_axi_awvalid),
    .m07_axi_awready(m07_axi_awready),
    .m07_axi_awaddr(m07_axi_awaddr),
    .m07_axi_awlen(m07_axi_awlen),
    .m07_axi_wvalid(m07_axi_wvalid),
    .m07_axi_wready(m07_axi_wready),
    .m07_axi_wdata(m07_axi_wdata),
    .m07_axi_wstrb(m07_axi_wstrb),
    .m07_axi_wlast(m07_axi_wlast),
    .m07_axi_bvalid(m07_axi_bvalid),
    .m07_axi_bready(m07_axi_bready),
    .m07_axi_arvalid(m07_axi_arvalid),
    .m07_axi_arready(m07_axi_arready),
    .m07_axi_araddr(m07_axi_araddr),
    .m07_axi_arlen(m07_axi_arlen),
    .m07_axi_rvalid(m07_axi_rvalid),
    .m07_axi_rready(m07_axi_rready),
    .m07_axi_rdata(m07_axi_rdata),
    .m07_axi_rlast(m07_axi_rlast),
    .m08_axi_awvalid(m08_axi_awvalid),
    .m08_axi_awready(m08_axi_awready),
    .m08_axi_awaddr(m08_axi_awaddr),
    .m08_axi_awlen(m08_axi_awlen),
    .m08_axi_wvalid(m08_axi_wvalid),
    .m08_axi_wready(m08_axi_wready),
    .m08_axi_wdata(m08_axi_wdata),
    .m08_axi_wstrb(m08_axi_wstrb),
    .m08_axi_wlast(m08_axi_wlast),
    .m08_axi_bvalid(m08_axi_bvalid),
    .m08_axi_bready(m08_axi_bready),
    .m08_axi_arvalid(m08_axi_arvalid),
    .m08_axi_arready(m08_axi_arready),
    .m08_axi_araddr(m08_axi_araddr),
    .m08_axi_arlen(m08_axi_arlen),
    .m08_axi_rvalid(m08_axi_rvalid),
    .m08_axi_rready(m08_axi_rready),
    .m08_axi_rdata(m08_axi_rdata),
    .m08_axi_rlast(m08_axi_rlast),
    .m09_axi_awvalid(m09_axi_awvalid),
    .m09_axi_awready(m09_axi_awready),
    .m09_axi_awaddr(m09_axi_awaddr),
    .m09_axi_awlen(m09_axi_awlen),
    .m09_axi_wvalid(m09_axi_wvalid),
    .m09_axi_wready(m09_axi_wready),
    .m09_axi_wdata(m09_axi_wdata),
    .m09_axi_wstrb(m09_axi_wstrb),
    .m09_axi_wlast(m09_axi_wlast),
    .m09_axi_bvalid(m09_axi_bvalid),
    .m09_axi_bready(m09_axi_bready),
    .m09_axi_arvalid(m09_axi_arvalid),
    .m09_axi_arready(m09_axi_arready),
    .m09_axi_araddr(m09_axi_araddr),
    .m09_axi_arlen(m09_axi_arlen),
    .m09_axi_rvalid(m09_axi_rvalid),
    .m09_axi_rready(m09_axi_rready),
    .m09_axi_rdata(m09_axi_rdata),
    .m09_axi_rlast(m09_axi_rlast),
    .m10_axi_awvalid(m10_axi_awvalid),
    .m10_axi_awready(m10_axi_awready),
    .m10_axi_awaddr(m10_axi_awaddr),
    .m10_axi_awlen(m10_axi_awlen),
    .m10_axi_wvalid(m10_axi_wvalid),
    .m10_axi_wready(m10_axi_wready),
    .m10_axi_wdata(m10_axi_wdata),
    .m10_axi_wstrb(m10_axi_wstrb),
    .m10_axi_wlast(m10_axi_wlast),
    .m10_axi_bvalid(m10_axi_bvalid),
    .m10_axi_bready(m10_axi_bready),
    .m10_axi_arvalid(m10_axi_arvalid),
    .m10_axi_arready(m10_axi_arready),
    .m10_axi_araddr(m10_axi_araddr),
    .m10_axi_arlen(m10_axi_arlen),
    .m10_axi_rvalid(m10_axi_rvalid),
    .m10_axi_rready(m10_axi_rready),
    .m10_axi_rdata(m10_axi_rdata),
    .m10_axi_rlast(m10_axi_rlast),
    .m11_axi_awvalid(m11_axi_awvalid),
    .m11_axi_awready(m11_axi_awready),
    .m11_axi_awaddr(m11_axi_awaddr),
    .m11_axi_awlen(m11_axi_awlen),
    .m11_axi_wvalid(m11_axi_wvalid),
    .m11_axi_wready(m11_axi_wready),
    .m11_axi_wdata(m11_axi_wdata),
    .m11_axi_wstrb(m11_axi_wstrb),
    .m11_axi_wlast(m11_axi_wlast),
    .m11_axi_bvalid(m11_axi_bvalid),
    .m11_axi_bready(m11_axi_bready),
    .m11_axi_arvalid(m11_axi_arvalid),
    .m11_axi_arready(m11_axi_arready),
    .m11_axi_araddr(m11_axi_araddr),
    .m11_axi_arlen(m11_axi_arlen),
    .m11_axi_rvalid(m11_axi_rvalid),
    .m11_axi_rready(m11_axi_rready),
    .m11_axi_rdata(m11_axi_rdata),
    .m11_axi_rlast(m11_axi_rlast),
    .m12_axi_awvalid(m12_axi_awvalid),
    .m12_axi_awready(m12_axi_awready),
    .m12_axi_awaddr(m12_axi_awaddr),
    .m12_axi_awlen(m12_axi_awlen),
    .m12_axi_wvalid(m12_axi_wvalid),
    .m12_axi_wready(m12_axi_wready),
    .m12_axi_wdata(m12_axi_wdata),
    .m12_axi_wstrb(m12_axi_wstrb),
    .m12_axi_wlast(m12_axi_wlast),
    .m12_axi_bvalid(m12_axi_bvalid),
    .m12_axi_bready(m12_axi_bready),
    .m12_axi_arvalid(m12_axi_arvalid),
    .m12_axi_arready(m12_axi_arready),
    .m12_axi_araddr(m12_axi_araddr),
    .m12_axi_arlen(m12_axi_arlen),
    .m12_axi_rvalid(m12_axi_rvalid),
    .m12_axi_rready(m12_axi_rready),
    .m12_axi_rdata(m12_axi_rdata),
    .m12_axi_rlast(m12_axi_rlast),
    .m13_axi_awvalid(m13_axi_awvalid),
    .m13_axi_awready(m13_axi_awready),
    .m13_axi_awaddr(m13_axi_awaddr),
    .m13_axi_awlen(m13_axi_awlen),
    .m13_axi_wvalid(m13_axi_wvalid),
    .m13_axi_wready(m13_axi_wready),
    .m13_axi_wdata(m13_axi_wdata),
    .m13_axi_wstrb(m13_axi_wstrb),
    .m13_axi_wlast(m13_axi_wlast),
    .m13_axi_bvalid(m13_axi_bvalid),
    .m13_axi_bready(m13_axi_bready),
    .m13_axi_arvalid(m13_axi_arvalid),
    .m13_axi_arready(m13_axi_arready),
    .m13_axi_araddr(m13_axi_araddr),
    .m13_axi_arlen(m13_axi_arlen),
    .m13_axi_rvalid(m13_axi_rvalid),
    .m13_axi_rready(m13_axi_rready),
    .m13_axi_rdata(m13_axi_rdata),
    .m13_axi_rlast(m13_axi_rlast),
    .m14_axi_awvalid(m14_axi_awvalid),
    .m14_axi_awready(m14_axi_awready),
    .m14_axi_awaddr(m14_axi_awaddr),
    .m14_axi_awlen(m14_axi_awlen),
    .m14_axi_wvalid(m14_axi_wvalid),
    .m14_axi_wready(m14_axi_wready),
    .m14_axi_wdata(m14_axi_wdata),
    .m14_axi_wstrb(m14_axi_wstrb),
    .m14_axi_wlast(m14_axi_wlast),
    .m14_axi_bvalid(m14_axi_bvalid),
    .m14_axi_bready(m14_axi_bready),
    .m14_axi_arvalid(m14_axi_arvalid),
    .m14_axi_arready(m14_axi_arready),
    .m14_axi_araddr(m14_axi_araddr),
    .m14_axi_arlen(m14_axi_arlen),
    .m14_axi_rvalid(m14_axi_rvalid),
    .m14_axi_rready(m14_axi_rready),
    .m14_axi_rdata(m14_axi_rdata),
    .m14_axi_rlast(m14_axi_rlast),
    .m15_axi_awvalid(m15_axi_awvalid),
    .m15_axi_awready(m15_axi_awready),
    .m15_axi_awaddr(m15_axi_awaddr),
    .m15_axi_awlen(m15_axi_awlen),
    .m15_axi_wvalid(m15_axi_wvalid),
    .m15_axi_wready(m15_axi_wready),
    .m15_axi_wdata(m15_axi_wdata),
    .m15_axi_wstrb(m15_axi_wstrb),
    .m15_axi_wlast(m15_axi_wlast),
    .m15_axi_bvalid(m15_axi_bvalid),
    .m15_axi_bready(m15_axi_bready),
    .m15_axi_arvalid(m15_axi_arvalid),
    .m15_axi_arready(m15_axi_arready),
    .m15_axi_araddr(m15_axi_araddr),
    .m15_axi_arlen(m15_axi_arlen),
    .m15_axi_rvalid(m15_axi_rvalid),
    .m15_axi_rready(m15_axi_rready),
    .m15_axi_rdata(m15_axi_rdata),
    .m15_axi_rlast(m15_axi_rlast),
    .m16_axi_awvalid(m16_axi_awvalid),
    .m16_axi_awready(m16_axi_awready),
    .m16_axi_awaddr(m16_axi_awaddr),
    .m16_axi_awlen(m16_axi_awlen),
    .m16_axi_wvalid(m16_axi_wvalid),
    .m16_axi_wready(m16_axi_wready),
    .m16_axi_wdata(m16_axi_wdata),
    .m16_axi_wstrb(m16_axi_wstrb),
    .m16_axi_wlast(m16_axi_wlast),
    .m16_axi_bvalid(m16_axi_bvalid),
    .m16_axi_bready(m16_axi_bready),
    .m16_axi_arvalid(m16_axi_arvalid),
    .m16_axi_arready(m16_axi_arready),
    .m16_axi_araddr(m16_axi_araddr),
    .m16_axi_arlen(m16_axi_arlen),
    .m16_axi_rvalid(m16_axi_rvalid),
    .m16_axi_rready(m16_axi_rready),
    .m16_axi_rdata(m16_axi_rdata),
    .m16_axi_rlast(m16_axi_rlast),
    .m17_axi_awvalid(m17_axi_awvalid),
    .m17_axi_awready(m17_axi_awready),
    .m17_axi_awaddr(m17_axi_awaddr),
    .m17_axi_awlen(m17_axi_awlen),
    .m17_axi_wvalid(m17_axi_wvalid),
    .m17_axi_wready(m17_axi_wready),
    .m17_axi_wdata(m17_axi_wdata),
    .m17_axi_wstrb(m17_axi_wstrb),
    .m17_axi_wlast(m17_axi_wlast),
    .m17_axi_bvalid(m17_axi_bvalid),
    .m17_axi_bready(m17_axi_bready),
    .m17_axi_arvalid(m17_axi_arvalid),
    .m17_axi_arready(m17_axi_arready),
    .m17_axi_araddr(m17_axi_araddr),
    .m17_axi_arlen(m17_axi_arlen),
    .m17_axi_rvalid(m17_axi_rvalid),
    .m17_axi_rready(m17_axi_rready),
    .m17_axi_rdata(m17_axi_rdata),
    .m17_axi_rlast(m17_axi_rlast),
    .m18_axi_awvalid(m18_axi_awvalid),
    .m18_axi_awready(m18_axi_awready),
    .m18_axi_awaddr(m18_axi_awaddr),
    .m18_axi_awlen(m18_axi_awlen),
    .m18_axi_wvalid(m18_axi_wvalid),
    .m18_axi_wready(m18_axi_wready),
    .m18_axi_wdata(m18_axi_wdata),
    .m18_axi_wstrb(m18_axi_wstrb),
    .m18_axi_wlast(m18_axi_wlast),
    .m18_axi_bvalid(m18_axi_bvalid),
    .m18_axi_bready(m18_axi_bready),
    .m18_axi_arvalid(m18_axi_arvalid),
    .m18_axi_arready(m18_axi_arready),
    .m18_axi_araddr(m18_axi_araddr),
    .m18_axi_arlen(m18_axi_arlen),
    .m18_axi_rvalid(m18_axi_rvalid),
    .m18_axi_rready(m18_axi_rready),
    .m18_axi_rdata(m18_axi_rdata),
    .m18_axi_rlast(m18_axi_rlast),
    .m19_axi_awvalid(m19_axi_awvalid),
    .m19_axi_awready(m19_axi_awready),
    .m19_axi_awaddr(m19_axi_awaddr),
    .m19_axi_awlen(m19_axi_awlen),
    .m19_axi_wvalid(m19_axi_wvalid),
    .m19_axi_wready(m19_axi_wready),
    .m19_axi_wdata(m19_axi_wdata),
    .m19_axi_wstrb(m19_axi_wstrb),
    .m19_axi_wlast(m19_axi_wlast),
    .m19_axi_bvalid(m19_axi_bvalid),
    .m19_axi_bready(m19_axi_bready),
    .m19_axi_arvalid(m19_axi_arvalid),
    .m19_axi_arready(m19_axi_arready),
    .m19_axi_araddr(m19_axi_araddr),
    .m19_axi_arlen(m19_axi_arlen),
    .m19_axi_rvalid(m19_axi_rvalid),
    .m19_axi_rready(m19_axi_rready),
    .m19_axi_rdata(m19_axi_rdata),
    .m19_axi_rlast(m19_axi_rlast),
    .m20_axi_awvalid(m20_axi_awvalid),
    .m20_axi_awready(m20_axi_awready),
    .m20_axi_awaddr(m20_axi_awaddr),
    .m20_axi_awlen(m20_axi_awlen),
    .m20_axi_wvalid(m20_axi_wvalid),
    .m20_axi_wready(m20_axi_wready),
    .m20_axi_wdata(m20_axi_wdata),
    .m20_axi_wstrb(m20_axi_wstrb),
    .m20_axi_wlast(m20_axi_wlast),
    .m20_axi_bvalid(m20_axi_bvalid),
    .m20_axi_bready(m20_axi_bready),
    .m20_axi_arvalid(m20_axi_arvalid),
    .m20_axi_arready(m20_axi_arready),
    .m20_axi_araddr(m20_axi_araddr),
    .m20_axi_arlen(m20_axi_arlen),
    .m20_axi_rvalid(m20_axi_rvalid),
    .m20_axi_rready(m20_axi_rready),
    .m20_axi_rdata(m20_axi_rdata),
    .m20_axi_rlast(m20_axi_rlast),
    .m21_axi_awvalid(m21_axi_awvalid),
    .m21_axi_awready(m21_axi_awready),
    .m21_axi_awaddr(m21_axi_awaddr),
    .m21_axi_awlen(m21_axi_awlen),
    .m21_axi_wvalid(m21_axi_wvalid),
    .m21_axi_wready(m21_axi_wready),
    .m21_axi_wdata(m21_axi_wdata),
    .m21_axi_wstrb(m21_axi_wstrb),
    .m21_axi_wlast(m21_axi_wlast),
    .m21_axi_bvalid(m21_axi_bvalid),
    .m21_axi_bready(m21_axi_bready),
    .m21_axi_arvalid(m21_axi_arvalid),
    .m21_axi_arready(m21_axi_arready),
    .m21_axi_araddr(m21_axi_araddr),
    .m21_axi_arlen(m21_axi_arlen),
    .m21_axi_rvalid(m21_axi_rvalid),
    .m21_axi_rready(m21_axi_rready),
    .m21_axi_rdata(m21_axi_rdata),
    .m21_axi_rlast(m21_axi_rlast),
    .m22_axi_awvalid(m22_axi_awvalid),
    .m22_axi_awready(m22_axi_awready),
    .m22_axi_awaddr(m22_axi_awaddr),
    .m22_axi_awlen(m22_axi_awlen),
    .m22_axi_wvalid(m22_axi_wvalid),
    .m22_axi_wready(m22_axi_wready),
    .m22_axi_wdata(m22_axi_wdata),
    .m22_axi_wstrb(m22_axi_wstrb),
    .m22_axi_wlast(m22_axi_wlast),
    .m22_axi_bvalid(m22_axi_bvalid),
    .m22_axi_bready(m22_axi_bready),
    .m22_axi_arvalid(m22_axi_arvalid),
    .m22_axi_arready(m22_axi_arready),
    .m22_axi_araddr(m22_axi_araddr),
    .m22_axi_arlen(m22_axi_arlen),
    .m22_axi_rvalid(m22_axi_rvalid),
    .m22_axi_rready(m22_axi_rready),
    .m22_axi_rdata(m22_axi_rdata),
    .m22_axi_rlast(m22_axi_rlast),
    .m23_axi_awvalid(m23_axi_awvalid),
    .m23_axi_awready(m23_axi_awready),
    .m23_axi_awaddr(m23_axi_awaddr),
    .m23_axi_awlen(m23_axi_awlen),
    .m23_axi_wvalid(m23_axi_wvalid),
    .m23_axi_wready(m23_axi_wready),
    .m23_axi_wdata(m23_axi_wdata),
    .m23_axi_wstrb(m23_axi_wstrb),
    .m23_axi_wlast(m23_axi_wlast),
    .m23_axi_bvalid(m23_axi_bvalid),
    .m23_axi_bready(m23_axi_bready),
    .m23_axi_arvalid(m23_axi_arvalid),
    .m23_axi_arready(m23_axi_arready),
    .m23_axi_araddr(m23_axi_araddr),
    .m23_axi_arlen(m23_axi_arlen),
    .m23_axi_rvalid(m23_axi_rvalid),
    .m23_axi_rready(m23_axi_rready),
    .m23_axi_rdata(m23_axi_rdata),
    .m23_axi_rlast(m23_axi_rlast),
    .m24_axi_awvalid(m24_axi_awvalid),
    .m24_axi_awready(m24_axi_awready),
    .m24_axi_awaddr(m24_axi_awaddr),
    .m24_axi_awlen(m24_axi_awlen),
    .m24_axi_wvalid(m24_axi_wvalid),
    .m24_axi_wready(m24_axi_wready),
    .m24_axi_wdata(m24_axi_wdata),
    .m24_axi_wstrb(m24_axi_wstrb),
    .m24_axi_wlast(m24_axi_wlast),
    .m24_axi_bvalid(m24_axi_bvalid),
    .m24_axi_bready(m24_axi_bready),
    .m24_axi_arvalid(m24_axi_arvalid),
    .m24_axi_arready(m24_axi_arready),
    .m24_axi_araddr(m24_axi_araddr),
    .m24_axi_arlen(m24_axi_arlen),
    .m24_axi_rvalid(m24_axi_rvalid),
    .m24_axi_rready(m24_axi_rready),
    .m24_axi_rdata(m24_axi_rdata),
    .m24_axi_rlast(m24_axi_rlast),
    .m25_axi_awvalid(m25_axi_awvalid),
    .m25_axi_awready(m25_axi_awready),
    .m25_axi_awaddr(m25_axi_awaddr),
    .m25_axi_awlen(m25_axi_awlen),
    .m25_axi_wvalid(m25_axi_wvalid),
    .m25_axi_wready(m25_axi_wready),
    .m25_axi_wdata(m25_axi_wdata),
    .m25_axi_wstrb(m25_axi_wstrb),
    .m25_axi_wlast(m25_axi_wlast),
    .m25_axi_bvalid(m25_axi_bvalid),
    .m25_axi_bready(m25_axi_bready),
    .m25_axi_arvalid(m25_axi_arvalid),
    .m25_axi_arready(m25_axi_arready),
    .m25_axi_araddr(m25_axi_araddr),
    .m25_axi_arlen(m25_axi_arlen),
    .m25_axi_rvalid(m25_axi_rvalid),
    .m25_axi_rready(m25_axi_rready),
    .m25_axi_rdata(m25_axi_rdata),
    .m25_axi_rlast(m25_axi_rlast),
    .m26_axi_awvalid(m26_axi_awvalid),
    .m26_axi_awready(m26_axi_awready),
    .m26_axi_awaddr(m26_axi_awaddr),
    .m26_axi_awlen(m26_axi_awlen),
    .m26_axi_wvalid(m26_axi_wvalid),
    .m26_axi_wready(m26_axi_wready),
    .m26_axi_wdata(m26_axi_wdata),
    .m26_axi_wstrb(m26_axi_wstrb),
    .m26_axi_wlast(m26_axi_wlast),
    .m26_axi_bvalid(m26_axi_bvalid),
    .m26_axi_bready(m26_axi_bready),
    .m26_axi_arvalid(m26_axi_arvalid),
    .m26_axi_arready(m26_axi_arready),
    .m26_axi_araddr(m26_axi_araddr),
    .m26_axi_arlen(m26_axi_arlen),
    .m26_axi_rvalid(m26_axi_rvalid),
    .m26_axi_rready(m26_axi_rready),
    .m26_axi_rdata(m26_axi_rdata),
    .m26_axi_rlast(m26_axi_rlast),
    .m27_axi_awvalid(m27_axi_awvalid),
    .m27_axi_awready(m27_axi_awready),
    .m27_axi_awaddr(m27_axi_awaddr),
    .m27_axi_awlen(m27_axi_awlen),
    .m27_axi_wvalid(m27_axi_wvalid),
    .m27_axi_wready(m27_axi_wready),
    .m27_axi_wdata(m27_axi_wdata),
    .m27_axi_wstrb(m27_axi_wstrb),
    .m27_axi_wlast(m27_axi_wlast),
    .m27_axi_bvalid(m27_axi_bvalid),
    .m27_axi_bready(m27_axi_bready),
    .m27_axi_arvalid(m27_axi_arvalid),
    .m27_axi_arready(m27_axi_arready),
    .m27_axi_araddr(m27_axi_araddr),
    .m27_axi_arlen(m27_axi_arlen),
    .m27_axi_rvalid(m27_axi_rvalid),
    .m27_axi_rready(m27_axi_rready),
    .m27_axi_rdata(m27_axi_rdata),
    .m27_axi_rlast(m27_axi_rlast),
    .m28_axi_awvalid(m28_axi_awvalid),
    .m28_axi_awready(m28_axi_awready),
    .m28_axi_awaddr(m28_axi_awaddr),
    .m28_axi_awlen(m28_axi_awlen),
    .m28_axi_wvalid(m28_axi_wvalid),
    .m28_axi_wready(m28_axi_wready),
    .m28_axi_wdata(m28_axi_wdata),
    .m28_axi_wstrb(m28_axi_wstrb),
    .m28_axi_wlast(m28_axi_wlast),
    .m28_axi_bvalid(m28_axi_bvalid),
    .m28_axi_bready(m28_axi_bready),
    .m28_axi_arvalid(m28_axi_arvalid),
    .m28_axi_arready(m28_axi_arready),
    .m28_axi_araddr(m28_axi_araddr),
    .m28_axi_arlen(m28_axi_arlen),
    .m28_axi_rvalid(m28_axi_rvalid),
    .m28_axi_rready(m28_axi_rready),
    .m28_axi_rdata(m28_axi_rdata),
    .m28_axi_rlast(m28_axi_rlast),
    .m29_axi_awvalid(m29_axi_awvalid),
    .m29_axi_awready(m29_axi_awready),
    .m29_axi_awaddr(m29_axi_awaddr),
    .m29_axi_awlen(m29_axi_awlen),
    .m29_axi_wvalid(m29_axi_wvalid),
    .m29_axi_wready(m29_axi_wready),
    .m29_axi_wdata(m29_axi_wdata),
    .m29_axi_wstrb(m29_axi_wstrb),
    .m29_axi_wlast(m29_axi_wlast),
    .m29_axi_bvalid(m29_axi_bvalid),
    .m29_axi_bready(m29_axi_bready),
    .m29_axi_arvalid(m29_axi_arvalid),
    .m29_axi_arready(m29_axi_arready),
    .m29_axi_araddr(m29_axi_araddr),
    .m29_axi_arlen(m29_axi_arlen),
    .m29_axi_rvalid(m29_axi_rvalid),
    .m29_axi_rready(m29_axi_rready),
    .m29_axi_rdata(m29_axi_rdata),
    .m29_axi_rlast(m29_axi_rlast),
    .m30_axi_awvalid(m30_axi_awvalid),
    .m30_axi_awready(m30_axi_awready),
    .m30_axi_awaddr(m30_axi_awaddr),
    .m30_axi_awlen(m30_axi_awlen),
    .m30_axi_wvalid(m30_axi_wvalid),
    .m30_axi_wready(m30_axi_wready),
    .m30_axi_wdata(m30_axi_wdata),
    .m30_axi_wstrb(m30_axi_wstrb),
    .m30_axi_wlast(m30_axi_wlast),
    .m30_axi_bvalid(m30_axi_bvalid),
    .m30_axi_bready(m30_axi_bready),
    .m30_axi_arvalid(m30_axi_arvalid),
    .m30_axi_arready(m30_axi_arready),
    .m30_axi_araddr(m30_axi_araddr),
    .m30_axi_arlen(m30_axi_arlen),
    .m30_axi_rvalid(m30_axi_rvalid),
    .m30_axi_rready(m30_axi_rready),
    .m30_axi_rdata(m30_axi_rdata),
    .m30_axi_rlast(m30_axi_rlast),
    .m31_axi_awvalid(m31_axi_awvalid),
    .m31_axi_awready(m31_axi_awready),
    .m31_axi_awaddr(m31_axi_awaddr),
    .m31_axi_awlen(m31_axi_awlen),
    .m31_axi_wvalid(m31_axi_wvalid),
    .m31_axi_wready(m31_axi_wready),
    .m31_axi_wdata(m31_axi_wdata),
    .m31_axi_wstrb(m31_axi_wstrb),
    .m31_axi_wlast(m31_axi_wlast),
    .m31_axi_bvalid(m31_axi_bvalid),
    .m31_axi_bready(m31_axi_bready),
    .m31_axi_arvalid(m31_axi_arvalid),
    .m31_axi_arready(m31_axi_arready),
    .m31_axi_araddr(m31_axi_araddr),
    .m31_axi_arlen(m31_axi_arlen),
    .m31_axi_rvalid(m31_axi_rvalid),
    .m31_axi_rready(m31_axi_rready),
    .m31_axi_rdata(m31_axi_rdata),
    .m31_axi_rlast(m31_axi_rlast)
  );


  initial begin
    areset = 1'b1;
  end


endmodule



module control_s_axi_32 #
(
  parameter C_S_AXI_ADDR_WIDTH = 11,
  parameter C_S_AXI_DATA_WIDTH = 32
)
(
  input aclk,
  input areset,
  input aclk_en,
  input [C_S_AXI_ADDR_WIDTH-1:0] awaddr,
  input awvalid,
  output awready,
  input [C_S_AXI_DATA_WIDTH-1:0] wdata,
  input [C_S_AXI_DATA_WIDTH/8-1:0] wstrb,
  input wvalid,
  output wready,
  output [2-1:0] bresp,
  output bvalid,
  input bready,
  input [C_S_AXI_ADDR_WIDTH-1:0] araddr,
  input arvalid,
  output arready,
  output [C_S_AXI_DATA_WIDTH-1:0] rdata,
  output [2-1:0] rresp,
  output rvalid,
  input rready,
  output interrupt,
  output ap_start,
  input ap_done,
  input ap_ready,
  input ap_idle,
  output [32-1:0] in_s0,
  output [32-1:0] in_s1,
  output [32-1:0] in_s2,
  output [32-1:0] in_s3,
  output [32-1:0] in_s4,
  output [32-1:0] in_s5,
  output [32-1:0] in_s6,
  output [32-1:0] in_s7,
  output [32-1:0] in_s8,
  output [32-1:0] in_s9,
  output [32-1:0] in_s10,
  output [32-1:0] in_s11,
  output [32-1:0] in_s12,
  output [32-1:0] in_s13,
  output [32-1:0] in_s14,
  output [32-1:0] in_s15,
  output [32-1:0] in_s16,
  output [32-1:0] in_s17,
  output [32-1:0] in_s18,
  output [32-1:0] in_s19,
  output [32-1:0] in_s20,
  output [32-1:0] in_s21,
  output [32-1:0] in_s22,
  output [32-1:0] in_s23,
  output [32-1:0] in_s24,
  output [32-1:0] in_s25,
  output [32-1:0] in_s26,
  output [32-1:0] in_s27,
  output [32-1:0] in_s28,
  output [32-1:0] in_s29,
  output [32-1:0] in_s30,
  output [32-1:0] in_s31,
  output [32-1:0] out_s0,
  output [32-1:0] out_s1,
  output [32-1:0] out_s2,
  output [32-1:0] out_s3,
  output [32-1:0] out_s4,
  output [32-1:0] out_s5,
  output [32-1:0] out_s6,
  output [32-1:0] out_s7,
  output [32-1:0] out_s8,
  output [32-1:0] out_s9,
  output [32-1:0] out_s10,
  output [32-1:0] out_s11,
  output [32-1:0] out_s12,
  output [32-1:0] out_s13,
  output [32-1:0] out_s14,
  output [32-1:0] out_s15,
  output [32-1:0] out_s16,
  output [32-1:0] out_s17,
  output [32-1:0] out_s18,
  output [32-1:0] out_s19,
  output [32-1:0] out_s20,
  output [32-1:0] out_s21,
  output [32-1:0] out_s22,
  output [32-1:0] out_s23,
  output [32-1:0] out_s24,
  output [32-1:0] out_s25,
  output [32-1:0] out_s26,
  output [32-1:0] out_s27,
  output [32-1:0] out_s28,
  output [32-1:0] out_s29,
  output [32-1:0] out_s30,
  output [32-1:0] out_s31,
  output [64-1:0] in0,
  output [64-1:0] in1,
  output [64-1:0] in2,
  output [64-1:0] in3,
  output [64-1:0] in4,
  output [64-1:0] in5,
  output [64-1:0] in6,
  output [64-1:0] in7,
  output [64-1:0] in8,
  output [64-1:0] in9,
  output [64-1:0] in10,
  output [64-1:0] in11,
  output [64-1:0] in12,
  output [64-1:0] in13,
  output [64-1:0] in14,
  output [64-1:0] in15,
  output [64-1:0] in16,
  output [64-1:0] in17,
  output [64-1:0] in18,
  output [64-1:0] in19,
  output [64-1:0] in20,
  output [64-1:0] in21,
  output [64-1:0] in22,
  output [64-1:0] in23,
  output [64-1:0] in24,
  output [64-1:0] in25,
  output [64-1:0] in26,
  output [64-1:0] in27,
  output [64-1:0] in28,
  output [64-1:0] in29,
  output [64-1:0] in30,
  output [64-1:0] in31,
  output [64-1:0] out0,
  output [64-1:0] out1,
  output [64-1:0] out2,
  output [64-1:0] out3,
  output [64-1:0] out4,
  output [64-1:0] out5,
  output [64-1:0] out6,
  output [64-1:0] out7,
  output [64-1:0] out8,
  output [64-1:0] out9,
  output [64-1:0] out10,
  output [64-1:0] out11,
  output [64-1:0] out12,
  output [64-1:0] out13,
  output [64-1:0] out14,
  output [64-1:0] out15,
  output [64-1:0] out16,
  output [64-1:0] out17,
  output [64-1:0] out18,
  output [64-1:0] out19,
  output [64-1:0] out20,
  output [64-1:0] out21,
  output [64-1:0] out22,
  output [64-1:0] out23,
  output [64-1:0] out24,
  output [64-1:0] out25,
  output [64-1:0] out26,
  output [64-1:0] out27,
  output [64-1:0] out28,
  output [64-1:0] out29,
  output [64-1:0] out30,
  output [64-1:0] out31
);

  localparam ADDR_AP_CTRL = 11'h0;
  localparam ADDR_GIE = 11'h4;
  localparam ADDR_IER = 11'h8;
  localparam ADDR_ISR = 11'hc;
  localparam ADDR_IN_S0_DATA_0 = 11'h10;
  localparam ADDR_IN_S0_CTRL = 11'h14;
  localparam ADDR_IN_S1_DATA_0 = 11'h18;
  localparam ADDR_IN_S1_CTRL = 11'h1c;
  localparam ADDR_IN_S2_DATA_0 = 11'h20;
  localparam ADDR_IN_S2_CTRL = 11'h24;
  localparam ADDR_IN_S3_DATA_0 = 11'h28;
  localparam ADDR_IN_S3_CTRL = 11'h2c;
  localparam ADDR_IN_S4_DATA_0 = 11'h30;
  localparam ADDR_IN_S4_CTRL = 11'h34;
  localparam ADDR_IN_S5_DATA_0 = 11'h38;
  localparam ADDR_IN_S5_CTRL = 11'h3c;
  localparam ADDR_IN_S6_DATA_0 = 11'h40;
  localparam ADDR_IN_S6_CTRL = 11'h44;
  localparam ADDR_IN_S7_DATA_0 = 11'h48;
  localparam ADDR_IN_S7_CTRL = 11'h4c;
  localparam ADDR_IN_S8_DATA_0 = 11'h50;
  localparam ADDR_IN_S8_CTRL = 11'h54;
  localparam ADDR_IN_S9_DATA_0 = 11'h58;
  localparam ADDR_IN_S9_CTRL = 11'h5c;
  localparam ADDR_IN_S10_DATA_0 = 11'h60;
  localparam ADDR_IN_S10_CTRL = 11'h64;
  localparam ADDR_IN_S11_DATA_0 = 11'h68;
  localparam ADDR_IN_S11_CTRL = 11'h6c;
  localparam ADDR_IN_S12_DATA_0 = 11'h70;
  localparam ADDR_IN_S12_CTRL = 11'h74;
  localparam ADDR_IN_S13_DATA_0 = 11'h78;
  localparam ADDR_IN_S13_CTRL = 11'h7c;
  localparam ADDR_IN_S14_DATA_0 = 11'h80;
  localparam ADDR_IN_S14_CTRL = 11'h84;
  localparam ADDR_IN_S15_DATA_0 = 11'h88;
  localparam ADDR_IN_S15_CTRL = 11'h8c;
  localparam ADDR_IN_S16_DATA_0 = 11'h90;
  localparam ADDR_IN_S16_CTRL = 11'h94;
  localparam ADDR_IN_S17_DATA_0 = 11'h98;
  localparam ADDR_IN_S17_CTRL = 11'h9c;
  localparam ADDR_IN_S18_DATA_0 = 11'ha0;
  localparam ADDR_IN_S18_CTRL = 11'ha4;
  localparam ADDR_IN_S19_DATA_0 = 11'ha8;
  localparam ADDR_IN_S19_CTRL = 11'hac;
  localparam ADDR_IN_S20_DATA_0 = 11'hb0;
  localparam ADDR_IN_S20_CTRL = 11'hb4;
  localparam ADDR_IN_S21_DATA_0 = 11'hb8;
  localparam ADDR_IN_S21_CTRL = 11'hbc;
  localparam ADDR_IN_S22_DATA_0 = 11'hc0;
  localparam ADDR_IN_S22_CTRL = 11'hc4;
  localparam ADDR_IN_S23_DATA_0 = 11'hc8;
  localparam ADDR_IN_S23_CTRL = 11'hcc;
  localparam ADDR_IN_S24_DATA_0 = 11'hd0;
  localparam ADDR_IN_S24_CTRL = 11'hd4;
  localparam ADDR_IN_S25_DATA_0 = 11'hd8;
  localparam ADDR_IN_S25_CTRL = 11'hdc;
  localparam ADDR_IN_S26_DATA_0 = 11'he0;
  localparam ADDR_IN_S26_CTRL = 11'he4;
  localparam ADDR_IN_S27_DATA_0 = 11'he8;
  localparam ADDR_IN_S27_CTRL = 11'hec;
  localparam ADDR_IN_S28_DATA_0 = 11'hf0;
  localparam ADDR_IN_S28_CTRL = 11'hf4;
  localparam ADDR_IN_S29_DATA_0 = 11'hf8;
  localparam ADDR_IN_S29_CTRL = 11'hfc;
  localparam ADDR_IN_S30_DATA_0 = 11'h100;
  localparam ADDR_IN_S30_CTRL = 11'h104;
  localparam ADDR_IN_S31_DATA_0 = 11'h108;
  localparam ADDR_IN_S31_CTRL = 11'h10c;
  localparam ADDR_OUT_S0_DATA_0 = 11'h110;
  localparam ADDR_OUT_S0_CTRL = 11'h114;
  localparam ADDR_OUT_S1_DATA_0 = 11'h118;
  localparam ADDR_OUT_S1_CTRL = 11'h11c;
  localparam ADDR_OUT_S2_DATA_0 = 11'h120;
  localparam ADDR_OUT_S2_CTRL = 11'h124;
  localparam ADDR_OUT_S3_DATA_0 = 11'h128;
  localparam ADDR_OUT_S3_CTRL = 11'h12c;
  localparam ADDR_OUT_S4_DATA_0 = 11'h130;
  localparam ADDR_OUT_S4_CTRL = 11'h134;
  localparam ADDR_OUT_S5_DATA_0 = 11'h138;
  localparam ADDR_OUT_S5_CTRL = 11'h13c;
  localparam ADDR_OUT_S6_DATA_0 = 11'h140;
  localparam ADDR_OUT_S6_CTRL = 11'h144;
  localparam ADDR_OUT_S7_DATA_0 = 11'h148;
  localparam ADDR_OUT_S7_CTRL = 11'h14c;
  localparam ADDR_OUT_S8_DATA_0 = 11'h150;
  localparam ADDR_OUT_S8_CTRL = 11'h154;
  localparam ADDR_OUT_S9_DATA_0 = 11'h158;
  localparam ADDR_OUT_S9_CTRL = 11'h15c;
  localparam ADDR_OUT_S10_DATA_0 = 11'h160;
  localparam ADDR_OUT_S10_CTRL = 11'h164;
  localparam ADDR_OUT_S11_DATA_0 = 11'h168;
  localparam ADDR_OUT_S11_CTRL = 11'h16c;
  localparam ADDR_OUT_S12_DATA_0 = 11'h170;
  localparam ADDR_OUT_S12_CTRL = 11'h174;
  localparam ADDR_OUT_S13_DATA_0 = 11'h178;
  localparam ADDR_OUT_S13_CTRL = 11'h17c;
  localparam ADDR_OUT_S14_DATA_0 = 11'h180;
  localparam ADDR_OUT_S14_CTRL = 11'h184;
  localparam ADDR_OUT_S15_DATA_0 = 11'h188;
  localparam ADDR_OUT_S15_CTRL = 11'h18c;
  localparam ADDR_OUT_S16_DATA_0 = 11'h190;
  localparam ADDR_OUT_S16_CTRL = 11'h194;
  localparam ADDR_OUT_S17_DATA_0 = 11'h198;
  localparam ADDR_OUT_S17_CTRL = 11'h19c;
  localparam ADDR_OUT_S18_DATA_0 = 11'h1a0;
  localparam ADDR_OUT_S18_CTRL = 11'h1a4;
  localparam ADDR_OUT_S19_DATA_0 = 11'h1a8;
  localparam ADDR_OUT_S19_CTRL = 11'h1ac;
  localparam ADDR_OUT_S20_DATA_0 = 11'h1b0;
  localparam ADDR_OUT_S20_CTRL = 11'h1b4;
  localparam ADDR_OUT_S21_DATA_0 = 11'h1b8;
  localparam ADDR_OUT_S21_CTRL = 11'h1bc;
  localparam ADDR_OUT_S22_DATA_0 = 11'h1c0;
  localparam ADDR_OUT_S22_CTRL = 11'h1c4;
  localparam ADDR_OUT_S23_DATA_0 = 11'h1c8;
  localparam ADDR_OUT_S23_CTRL = 11'h1cc;
  localparam ADDR_OUT_S24_DATA_0 = 11'h1d0;
  localparam ADDR_OUT_S24_CTRL = 11'h1d4;
  localparam ADDR_OUT_S25_DATA_0 = 11'h1d8;
  localparam ADDR_OUT_S25_CTRL = 11'h1dc;
  localparam ADDR_OUT_S26_DATA_0 = 11'h1e0;
  localparam ADDR_OUT_S26_CTRL = 11'h1e4;
  localparam ADDR_OUT_S27_DATA_0 = 11'h1e8;
  localparam ADDR_OUT_S27_CTRL = 11'h1ec;
  localparam ADDR_OUT_S28_DATA_0 = 11'h1f0;
  localparam ADDR_OUT_S28_CTRL = 11'h1f4;
  localparam ADDR_OUT_S29_DATA_0 = 11'h1f8;
  localparam ADDR_OUT_S29_CTRL = 11'h1fc;
  localparam ADDR_OUT_S30_DATA_0 = 11'h200;
  localparam ADDR_OUT_S30_CTRL = 11'h204;
  localparam ADDR_OUT_S31_DATA_0 = 11'h208;
  localparam ADDR_OUT_S31_CTRL = 11'h20c;
  localparam ADDR_IN0_DATA_0 = 11'h210;
  localparam ADDR_IN0_DATA_1 = 11'h214;
  localparam ADDR_IN0_CTRL = 11'h218;
  localparam ADDR_OUT0_DATA_0 = 11'h21c;
  localparam ADDR_OUT0_DATA_1 = 11'h220;
  localparam ADDR_OUT0_CTRL = 11'h224;
  localparam ADDR_IN1_DATA_0 = 11'h228;
  localparam ADDR_IN1_DATA_1 = 11'h22c;
  localparam ADDR_IN1_CTRL = 11'h230;
  localparam ADDR_OUT1_DATA_0 = 11'h234;
  localparam ADDR_OUT1_DATA_1 = 11'h238;
  localparam ADDR_OUT1_CTRL = 11'h23c;
  localparam ADDR_IN2_DATA_0 = 11'h240;
  localparam ADDR_IN2_DATA_1 = 11'h244;
  localparam ADDR_IN2_CTRL = 11'h248;
  localparam ADDR_OUT2_DATA_0 = 11'h24c;
  localparam ADDR_OUT2_DATA_1 = 11'h250;
  localparam ADDR_OUT2_CTRL = 11'h254;
  localparam ADDR_IN3_DATA_0 = 11'h258;
  localparam ADDR_IN3_DATA_1 = 11'h25c;
  localparam ADDR_IN3_CTRL = 11'h260;
  localparam ADDR_OUT3_DATA_0 = 11'h264;
  localparam ADDR_OUT3_DATA_1 = 11'h268;
  localparam ADDR_OUT3_CTRL = 11'h26c;
  localparam ADDR_IN4_DATA_0 = 11'h270;
  localparam ADDR_IN4_DATA_1 = 11'h274;
  localparam ADDR_IN4_CTRL = 11'h278;
  localparam ADDR_OUT4_DATA_0 = 11'h27c;
  localparam ADDR_OUT4_DATA_1 = 11'h280;
  localparam ADDR_OUT4_CTRL = 11'h284;
  localparam ADDR_IN5_DATA_0 = 11'h288;
  localparam ADDR_IN5_DATA_1 = 11'h28c;
  localparam ADDR_IN5_CTRL = 11'h290;
  localparam ADDR_OUT5_DATA_0 = 11'h294;
  localparam ADDR_OUT5_DATA_1 = 11'h298;
  localparam ADDR_OUT5_CTRL = 11'h29c;
  localparam ADDR_IN6_DATA_0 = 11'h2a0;
  localparam ADDR_IN6_DATA_1 = 11'h2a4;
  localparam ADDR_IN6_CTRL = 11'h2a8;
  localparam ADDR_OUT6_DATA_0 = 11'h2ac;
  localparam ADDR_OUT6_DATA_1 = 11'h2b0;
  localparam ADDR_OUT6_CTRL = 11'h2b4;
  localparam ADDR_IN7_DATA_0 = 11'h2b8;
  localparam ADDR_IN7_DATA_1 = 11'h2bc;
  localparam ADDR_IN7_CTRL = 11'h2c0;
  localparam ADDR_OUT7_DATA_0 = 11'h2c4;
  localparam ADDR_OUT7_DATA_1 = 11'h2c8;
  localparam ADDR_OUT7_CTRL = 11'h2cc;
  localparam ADDR_IN8_DATA_0 = 11'h2d0;
  localparam ADDR_IN8_DATA_1 = 11'h2d4;
  localparam ADDR_IN8_CTRL = 11'h2d8;
  localparam ADDR_OUT8_DATA_0 = 11'h2dc;
  localparam ADDR_OUT8_DATA_1 = 11'h2e0;
  localparam ADDR_OUT8_CTRL = 11'h2e4;
  localparam ADDR_IN9_DATA_0 = 11'h2e8;
  localparam ADDR_IN9_DATA_1 = 11'h2ec;
  localparam ADDR_IN9_CTRL = 11'h2f0;
  localparam ADDR_OUT9_DATA_0 = 11'h2f4;
  localparam ADDR_OUT9_DATA_1 = 11'h2f8;
  localparam ADDR_OUT9_CTRL = 11'h2fc;
  localparam ADDR_IN10_DATA_0 = 11'h300;
  localparam ADDR_IN10_DATA_1 = 11'h304;
  localparam ADDR_IN10_CTRL = 11'h308;
  localparam ADDR_OUT10_DATA_0 = 11'h30c;
  localparam ADDR_OUT10_DATA_1 = 11'h310;
  localparam ADDR_OUT10_CTRL = 11'h314;
  localparam ADDR_IN11_DATA_0 = 11'h318;
  localparam ADDR_IN11_DATA_1 = 11'h31c;
  localparam ADDR_IN11_CTRL = 11'h320;
  localparam ADDR_OUT11_DATA_0 = 11'h324;
  localparam ADDR_OUT11_DATA_1 = 11'h328;
  localparam ADDR_OUT11_CTRL = 11'h32c;
  localparam ADDR_IN12_DATA_0 = 11'h330;
  localparam ADDR_IN12_DATA_1 = 11'h334;
  localparam ADDR_IN12_CTRL = 11'h338;
  localparam ADDR_OUT12_DATA_0 = 11'h33c;
  localparam ADDR_OUT12_DATA_1 = 11'h340;
  localparam ADDR_OUT12_CTRL = 11'h344;
  localparam ADDR_IN13_DATA_0 = 11'h348;
  localparam ADDR_IN13_DATA_1 = 11'h34c;
  localparam ADDR_IN13_CTRL = 11'h350;
  localparam ADDR_OUT13_DATA_0 = 11'h354;
  localparam ADDR_OUT13_DATA_1 = 11'h358;
  localparam ADDR_OUT13_CTRL = 11'h35c;
  localparam ADDR_IN14_DATA_0 = 11'h360;
  localparam ADDR_IN14_DATA_1 = 11'h364;
  localparam ADDR_IN14_CTRL = 11'h368;
  localparam ADDR_OUT14_DATA_0 = 11'h36c;
  localparam ADDR_OUT14_DATA_1 = 11'h370;
  localparam ADDR_OUT14_CTRL = 11'h374;
  localparam ADDR_IN15_DATA_0 = 11'h378;
  localparam ADDR_IN15_DATA_1 = 11'h37c;
  localparam ADDR_IN15_CTRL = 11'h380;
  localparam ADDR_OUT15_DATA_0 = 11'h384;
  localparam ADDR_OUT15_DATA_1 = 11'h388;
  localparam ADDR_OUT15_CTRL = 11'h38c;
  localparam ADDR_IN16_DATA_0 = 11'h390;
  localparam ADDR_IN16_DATA_1 = 11'h394;
  localparam ADDR_IN16_CTRL = 11'h398;
  localparam ADDR_OUT16_DATA_0 = 11'h39c;
  localparam ADDR_OUT16_DATA_1 = 11'h3a0;
  localparam ADDR_OUT16_CTRL = 11'h3a4;
  localparam ADDR_IN17_DATA_0 = 11'h3a8;
  localparam ADDR_IN17_DATA_1 = 11'h3ac;
  localparam ADDR_IN17_CTRL = 11'h3b0;
  localparam ADDR_OUT17_DATA_0 = 11'h3b4;
  localparam ADDR_OUT17_DATA_1 = 11'h3b8;
  localparam ADDR_OUT17_CTRL = 11'h3bc;
  localparam ADDR_IN18_DATA_0 = 11'h3c0;
  localparam ADDR_IN18_DATA_1 = 11'h3c4;
  localparam ADDR_IN18_CTRL = 11'h3c8;
  localparam ADDR_OUT18_DATA_0 = 11'h3cc;
  localparam ADDR_OUT18_DATA_1 = 11'h3d0;
  localparam ADDR_OUT18_CTRL = 11'h3d4;
  localparam ADDR_IN19_DATA_0 = 11'h3d8;
  localparam ADDR_IN19_DATA_1 = 11'h3dc;
  localparam ADDR_IN19_CTRL = 11'h3e0;
  localparam ADDR_OUT19_DATA_0 = 11'h3e4;
  localparam ADDR_OUT19_DATA_1 = 11'h3e8;
  localparam ADDR_OUT19_CTRL = 11'h3ec;
  localparam ADDR_IN20_DATA_0 = 11'h3f0;
  localparam ADDR_IN20_DATA_1 = 11'h3f4;
  localparam ADDR_IN20_CTRL = 11'h3f8;
  localparam ADDR_OUT20_DATA_0 = 11'h3fc;
  localparam ADDR_OUT20_DATA_1 = 11'h400;
  localparam ADDR_OUT20_CTRL = 11'h404;
  localparam ADDR_IN21_DATA_0 = 11'h408;
  localparam ADDR_IN21_DATA_1 = 11'h40c;
  localparam ADDR_IN21_CTRL = 11'h410;
  localparam ADDR_OUT21_DATA_0 = 11'h414;
  localparam ADDR_OUT21_DATA_1 = 11'h418;
  localparam ADDR_OUT21_CTRL = 11'h41c;
  localparam ADDR_IN22_DATA_0 = 11'h420;
  localparam ADDR_IN22_DATA_1 = 11'h424;
  localparam ADDR_IN22_CTRL = 11'h428;
  localparam ADDR_OUT22_DATA_0 = 11'h42c;
  localparam ADDR_OUT22_DATA_1 = 11'h430;
  localparam ADDR_OUT22_CTRL = 11'h434;
  localparam ADDR_IN23_DATA_0 = 11'h438;
  localparam ADDR_IN23_DATA_1 = 11'h43c;
  localparam ADDR_IN23_CTRL = 11'h440;
  localparam ADDR_OUT23_DATA_0 = 11'h444;
  localparam ADDR_OUT23_DATA_1 = 11'h448;
  localparam ADDR_OUT23_CTRL = 11'h44c;
  localparam ADDR_IN24_DATA_0 = 11'h450;
  localparam ADDR_IN24_DATA_1 = 11'h454;
  localparam ADDR_IN24_CTRL = 11'h458;
  localparam ADDR_OUT24_DATA_0 = 11'h45c;
  localparam ADDR_OUT24_DATA_1 = 11'h460;
  localparam ADDR_OUT24_CTRL = 11'h464;
  localparam ADDR_IN25_DATA_0 = 11'h468;
  localparam ADDR_IN25_DATA_1 = 11'h46c;
  localparam ADDR_IN25_CTRL = 11'h470;
  localparam ADDR_OUT25_DATA_0 = 11'h474;
  localparam ADDR_OUT25_DATA_1 = 11'h478;
  localparam ADDR_OUT25_CTRL = 11'h47c;
  localparam ADDR_IN26_DATA_0 = 11'h480;
  localparam ADDR_IN26_DATA_1 = 11'h484;
  localparam ADDR_IN26_CTRL = 11'h488;
  localparam ADDR_OUT26_DATA_0 = 11'h48c;
  localparam ADDR_OUT26_DATA_1 = 11'h490;
  localparam ADDR_OUT26_CTRL = 11'h494;
  localparam ADDR_IN27_DATA_0 = 11'h498;
  localparam ADDR_IN27_DATA_1 = 11'h49c;
  localparam ADDR_IN27_CTRL = 11'h4a0;
  localparam ADDR_OUT27_DATA_0 = 11'h4a4;
  localparam ADDR_OUT27_DATA_1 = 11'h4a8;
  localparam ADDR_OUT27_CTRL = 11'h4ac;
  localparam ADDR_IN28_DATA_0 = 11'h4b0;
  localparam ADDR_IN28_DATA_1 = 11'h4b4;
  localparam ADDR_IN28_CTRL = 11'h4b8;
  localparam ADDR_OUT28_DATA_0 = 11'h4bc;
  localparam ADDR_OUT28_DATA_1 = 11'h4c0;
  localparam ADDR_OUT28_CTRL = 11'h4c4;
  localparam ADDR_IN29_DATA_0 = 11'h4c8;
  localparam ADDR_IN29_DATA_1 = 11'h4cc;
  localparam ADDR_IN29_CTRL = 11'h4d0;
  localparam ADDR_OUT29_DATA_0 = 11'h4d4;
  localparam ADDR_OUT29_DATA_1 = 11'h4d8;
  localparam ADDR_OUT29_CTRL = 11'h4dc;
  localparam ADDR_IN30_DATA_0 = 11'h4e0;
  localparam ADDR_IN30_DATA_1 = 11'h4e4;
  localparam ADDR_IN30_CTRL = 11'h4e8;
  localparam ADDR_OUT30_DATA_0 = 11'h4ec;
  localparam ADDR_OUT30_DATA_1 = 11'h4f0;
  localparam ADDR_OUT30_CTRL = 11'h4f4;
  localparam ADDR_IN31_DATA_0 = 11'h4f8;
  localparam ADDR_IN31_DATA_1 = 11'h4fc;
  localparam ADDR_IN31_CTRL = 11'h500;
  localparam ADDR_OUT31_DATA_0 = 11'h504;
  localparam ADDR_OUT31_DATA_1 = 11'h508;
  localparam ADDR_OUT31_CTRL = 11'h50c;
  localparam WRIDLE = 2'd0;
  localparam WRDATA = 2'd1;
  localparam WRRESP = 2'd2;
  localparam WRRESET = 2'd3;
  localparam RDIDLE = 2'd0;
  localparam RDDATA = 2'd1;
  localparam RDRESET = 2'd2;
  localparam ADDR_BITS = 11;
  reg [2-1:0] wstate;
  reg [2-1:0] wnext;
  reg [ADDR_BITS-1:0] waddr;
  wire [32-1:0] wmask;
  wire aw_hs;
  wire w_hs;
  reg [2-1:0] rstate;
  reg [2-1:0] rnext;
  reg [32-1:0] rrdata;
  wire ar_hs;
  wire [ADDR_BITS-1:0] raddr;
  reg int_ap_idle;
  reg int_ap_ready;
  reg int_ap_done;
  reg int_ap_start;
  reg int_auto_restart;
  reg int_gie;
  reg [2-1:0] int_ier;
  reg [2-1:0] int_isr;
  reg [32-1:0] int_in_s0;
  reg [32-1:0] int_in_s1;
  reg [32-1:0] int_in_s2;
  reg [32-1:0] int_in_s3;
  reg [32-1:0] int_in_s4;
  reg [32-1:0] int_in_s5;
  reg [32-1:0] int_in_s6;
  reg [32-1:0] int_in_s7;
  reg [32-1:0] int_in_s8;
  reg [32-1:0] int_in_s9;
  reg [32-1:0] int_in_s10;
  reg [32-1:0] int_in_s11;
  reg [32-1:0] int_in_s12;
  reg [32-1:0] int_in_s13;
  reg [32-1:0] int_in_s14;
  reg [32-1:0] int_in_s15;
  reg [32-1:0] int_in_s16;
  reg [32-1:0] int_in_s17;
  reg [32-1:0] int_in_s18;
  reg [32-1:0] int_in_s19;
  reg [32-1:0] int_in_s20;
  reg [32-1:0] int_in_s21;
  reg [32-1:0] int_in_s22;
  reg [32-1:0] int_in_s23;
  reg [32-1:0] int_in_s24;
  reg [32-1:0] int_in_s25;
  reg [32-1:0] int_in_s26;
  reg [32-1:0] int_in_s27;
  reg [32-1:0] int_in_s28;
  reg [32-1:0] int_in_s29;
  reg [32-1:0] int_in_s30;
  reg [32-1:0] int_in_s31;
  reg [32-1:0] int_out_s0;
  reg [32-1:0] int_out_s1;
  reg [32-1:0] int_out_s2;
  reg [32-1:0] int_out_s3;
  reg [32-1:0] int_out_s4;
  reg [32-1:0] int_out_s5;
  reg [32-1:0] int_out_s6;
  reg [32-1:0] int_out_s7;
  reg [32-1:0] int_out_s8;
  reg [32-1:0] int_out_s9;
  reg [32-1:0] int_out_s10;
  reg [32-1:0] int_out_s11;
  reg [32-1:0] int_out_s12;
  reg [32-1:0] int_out_s13;
  reg [32-1:0] int_out_s14;
  reg [32-1:0] int_out_s15;
  reg [32-1:0] int_out_s16;
  reg [32-1:0] int_out_s17;
  reg [32-1:0] int_out_s18;
  reg [32-1:0] int_out_s19;
  reg [32-1:0] int_out_s20;
  reg [32-1:0] int_out_s21;
  reg [32-1:0] int_out_s22;
  reg [32-1:0] int_out_s23;
  reg [32-1:0] int_out_s24;
  reg [32-1:0] int_out_s25;
  reg [32-1:0] int_out_s26;
  reg [32-1:0] int_out_s27;
  reg [32-1:0] int_out_s28;
  reg [32-1:0] int_out_s29;
  reg [32-1:0] int_out_s30;
  reg [32-1:0] int_out_s31;
  reg [64-1:0] int_in0;
  reg [64-1:0] int_out0;
  reg [64-1:0] int_in1;
  reg [64-1:0] int_out1;
  reg [64-1:0] int_in2;
  reg [64-1:0] int_out2;
  reg [64-1:0] int_in3;
  reg [64-1:0] int_out3;
  reg [64-1:0] int_in4;
  reg [64-1:0] int_out4;
  reg [64-1:0] int_in5;
  reg [64-1:0] int_out5;
  reg [64-1:0] int_in6;
  reg [64-1:0] int_out6;
  reg [64-1:0] int_in7;
  reg [64-1:0] int_out7;
  reg [64-1:0] int_in8;
  reg [64-1:0] int_out8;
  reg [64-1:0] int_in9;
  reg [64-1:0] int_out9;
  reg [64-1:0] int_in10;
  reg [64-1:0] int_out10;
  reg [64-1:0] int_in11;
  reg [64-1:0] int_out11;
  reg [64-1:0] int_in12;
  reg [64-1:0] int_out12;
  reg [64-1:0] int_in13;
  reg [64-1:0] int_out13;
  reg [64-1:0] int_in14;
  reg [64-1:0] int_out14;
  reg [64-1:0] int_in15;
  reg [64-1:0] int_out15;
  reg [64-1:0] int_in16;
  reg [64-1:0] int_out16;
  reg [64-1:0] int_in17;
  reg [64-1:0] int_out17;
  reg [64-1:0] int_in18;
  reg [64-1:0] int_out18;
  reg [64-1:0] int_in19;
  reg [64-1:0] int_out19;
  reg [64-1:0] int_in20;
  reg [64-1:0] int_out20;
  reg [64-1:0] int_in21;
  reg [64-1:0] int_out21;
  reg [64-1:0] int_in22;
  reg [64-1:0] int_out22;
  reg [64-1:0] int_in23;
  reg [64-1:0] int_out23;
  reg [64-1:0] int_in24;
  reg [64-1:0] int_out24;
  reg [64-1:0] int_in25;
  reg [64-1:0] int_out25;
  reg [64-1:0] int_in26;
  reg [64-1:0] int_out26;
  reg [64-1:0] int_in27;
  reg [64-1:0] int_out27;
  reg [64-1:0] int_in28;
  reg [64-1:0] int_out28;
  reg [64-1:0] int_in29;
  reg [64-1:0] int_out29;
  reg [64-1:0] int_in30;
  reg [64-1:0] int_out30;
  reg [64-1:0] int_in31;
  reg [64-1:0] int_out31;
  assign awready = wstate == WRIDLE;
  assign wready = wstate == WRDATA;
  assign bresp = 2'b0;
  assign bvalid = wstate == WRRESP;
  assign wmask = { { 8{ wstrb[3] } }, { 8{ wstrb[2] } }, { 8{ wstrb[1] } }, { 8{ wstrb[0] } } };
  assign aw_hs = awvalid & awready;
  assign w_hs = wvalid & wready;

  always @(posedge aclk) begin
    if(areset) begin
      wstate <= WRRESET;
    end else begin
      if(aclk_en) begin
        wstate <= wnext;
      end 
    end
  end


  always @(*) begin
    case(wstate)
      WRIDLE: begin
        if(awvalid) begin
          wnext <= WRDATA;
        end else begin
          wnext <= WRIDLE;
        end
      end
      WRDATA: begin
        if(wvalid) begin
          wnext <= WRRESP;
        end else begin
          wnext <= WRDATA;
        end
      end
      WRRESP: begin
        if(bready) begin
          wnext <= WRIDLE;
        end else begin
          wnext <= WRRESP;
        end
      end
      default: begin
        wnext <= WRIDLE;
      end
    endcase
  end


  always @(posedge aclk) begin
    if(aclk_en) begin
      if(aw_hs) begin
        waddr <= awaddr[ADDR_BITS-1:0];
      end 
    end 
  end

  assign arready = rstate == RDIDLE;
  assign rdata = rrdata;
  assign rresp = 2'b0;
  assign rvalid = rstate == RDDATA;
  assign ar_hs = arvalid & arready;
  assign raddr = araddr[ADDR_BITS-1:0];

  always @(posedge aclk) begin
    if(areset) begin
      rstate <= RDRESET;
    end else begin
      if(aclk_en) begin
        rstate <= rnext;
      end 
    end
  end


  always @(*) begin
    case(rstate)
      RDIDLE: begin
        if(arvalid) begin
          rnext <= RDDATA;
        end else begin
          rnext <= RDIDLE;
        end
      end
      RDDATA: begin
        if(rready & rvalid) begin
          rnext <= RDIDLE;
        end else begin
          rnext <= RDDATA;
        end
      end
      default: begin
        rnext <= RDIDLE;
      end
    endcase
  end


  always @(posedge aclk) begin
    if(aclk_en) begin
      if(ar_hs) begin
        rrdata <= 1'b0;
        case(raddr)
          ADDR_AP_CTRL: begin
            rrdata[0] <= int_ap_start;
            rrdata[1] <= int_ap_done;
            rrdata[2] <= int_ap_idle;
            rrdata[3] <= int_ap_ready;
            rrdata[7] <= int_auto_restart;
          end
          ADDR_GIE: begin
            rrdata <= int_gie;
          end
          ADDR_IER: begin
            rrdata <= int_ier;
          end
          ADDR_ISR: begin
            rrdata <= int_isr;
          end
          ADDR_IN_S0_DATA_0: begin
            rrdata <= int_in_s0[31:0];
          end
          ADDR_IN_S1_DATA_0: begin
            rrdata <= int_in_s1[31:0];
          end
          ADDR_IN_S2_DATA_0: begin
            rrdata <= int_in_s2[31:0];
          end
          ADDR_IN_S3_DATA_0: begin
            rrdata <= int_in_s3[31:0];
          end
          ADDR_IN_S4_DATA_0: begin
            rrdata <= int_in_s4[31:0];
          end
          ADDR_IN_S5_DATA_0: begin
            rrdata <= int_in_s5[31:0];
          end
          ADDR_IN_S6_DATA_0: begin
            rrdata <= int_in_s6[31:0];
          end
          ADDR_IN_S7_DATA_0: begin
            rrdata <= int_in_s7[31:0];
          end
          ADDR_IN_S8_DATA_0: begin
            rrdata <= int_in_s8[31:0];
          end
          ADDR_IN_S9_DATA_0: begin
            rrdata <= int_in_s9[31:0];
          end
          ADDR_IN_S10_DATA_0: begin
            rrdata <= int_in_s10[31:0];
          end
          ADDR_IN_S11_DATA_0: begin
            rrdata <= int_in_s11[31:0];
          end
          ADDR_IN_S12_DATA_0: begin
            rrdata <= int_in_s12[31:0];
          end
          ADDR_IN_S13_DATA_0: begin
            rrdata <= int_in_s13[31:0];
          end
          ADDR_IN_S14_DATA_0: begin
            rrdata <= int_in_s14[31:0];
          end
          ADDR_IN_S15_DATA_0: begin
            rrdata <= int_in_s15[31:0];
          end
          ADDR_IN_S16_DATA_0: begin
            rrdata <= int_in_s16[31:0];
          end
          ADDR_IN_S17_DATA_0: begin
            rrdata <= int_in_s17[31:0];
          end
          ADDR_IN_S18_DATA_0: begin
            rrdata <= int_in_s18[31:0];
          end
          ADDR_IN_S19_DATA_0: begin
            rrdata <= int_in_s19[31:0];
          end
          ADDR_IN_S20_DATA_0: begin
            rrdata <= int_in_s20[31:0];
          end
          ADDR_IN_S21_DATA_0: begin
            rrdata <= int_in_s21[31:0];
          end
          ADDR_IN_S22_DATA_0: begin
            rrdata <= int_in_s22[31:0];
          end
          ADDR_IN_S23_DATA_0: begin
            rrdata <= int_in_s23[31:0];
          end
          ADDR_IN_S24_DATA_0: begin
            rrdata <= int_in_s24[31:0];
          end
          ADDR_IN_S25_DATA_0: begin
            rrdata <= int_in_s25[31:0];
          end
          ADDR_IN_S26_DATA_0: begin
            rrdata <= int_in_s26[31:0];
          end
          ADDR_IN_S27_DATA_0: begin
            rrdata <= int_in_s27[31:0];
          end
          ADDR_IN_S28_DATA_0: begin
            rrdata <= int_in_s28[31:0];
          end
          ADDR_IN_S29_DATA_0: begin
            rrdata <= int_in_s29[31:0];
          end
          ADDR_IN_S30_DATA_0: begin
            rrdata <= int_in_s30[31:0];
          end
          ADDR_IN_S31_DATA_0: begin
            rrdata <= int_in_s31[31:0];
          end
          ADDR_OUT_S0_DATA_0: begin
            rrdata <= int_out_s0[31:0];
          end
          ADDR_OUT_S1_DATA_0: begin
            rrdata <= int_out_s1[31:0];
          end
          ADDR_OUT_S2_DATA_0: begin
            rrdata <= int_out_s2[31:0];
          end
          ADDR_OUT_S3_DATA_0: begin
            rrdata <= int_out_s3[31:0];
          end
          ADDR_OUT_S4_DATA_0: begin
            rrdata <= int_out_s4[31:0];
          end
          ADDR_OUT_S5_DATA_0: begin
            rrdata <= int_out_s5[31:0];
          end
          ADDR_OUT_S6_DATA_0: begin
            rrdata <= int_out_s6[31:0];
          end
          ADDR_OUT_S7_DATA_0: begin
            rrdata <= int_out_s7[31:0];
          end
          ADDR_OUT_S8_DATA_0: begin
            rrdata <= int_out_s8[31:0];
          end
          ADDR_OUT_S9_DATA_0: begin
            rrdata <= int_out_s9[31:0];
          end
          ADDR_OUT_S10_DATA_0: begin
            rrdata <= int_out_s10[31:0];
          end
          ADDR_OUT_S11_DATA_0: begin
            rrdata <= int_out_s11[31:0];
          end
          ADDR_OUT_S12_DATA_0: begin
            rrdata <= int_out_s12[31:0];
          end
          ADDR_OUT_S13_DATA_0: begin
            rrdata <= int_out_s13[31:0];
          end
          ADDR_OUT_S14_DATA_0: begin
            rrdata <= int_out_s14[31:0];
          end
          ADDR_OUT_S15_DATA_0: begin
            rrdata <= int_out_s15[31:0];
          end
          ADDR_OUT_S16_DATA_0: begin
            rrdata <= int_out_s16[31:0];
          end
          ADDR_OUT_S17_DATA_0: begin
            rrdata <= int_out_s17[31:0];
          end
          ADDR_OUT_S18_DATA_0: begin
            rrdata <= int_out_s18[31:0];
          end
          ADDR_OUT_S19_DATA_0: begin
            rrdata <= int_out_s19[31:0];
          end
          ADDR_OUT_S20_DATA_0: begin
            rrdata <= int_out_s20[31:0];
          end
          ADDR_OUT_S21_DATA_0: begin
            rrdata <= int_out_s21[31:0];
          end
          ADDR_OUT_S22_DATA_0: begin
            rrdata <= int_out_s22[31:0];
          end
          ADDR_OUT_S23_DATA_0: begin
            rrdata <= int_out_s23[31:0];
          end
          ADDR_OUT_S24_DATA_0: begin
            rrdata <= int_out_s24[31:0];
          end
          ADDR_OUT_S25_DATA_0: begin
            rrdata <= int_out_s25[31:0];
          end
          ADDR_OUT_S26_DATA_0: begin
            rrdata <= int_out_s26[31:0];
          end
          ADDR_OUT_S27_DATA_0: begin
            rrdata <= int_out_s27[31:0];
          end
          ADDR_OUT_S28_DATA_0: begin
            rrdata <= int_out_s28[31:0];
          end
          ADDR_OUT_S29_DATA_0: begin
            rrdata <= int_out_s29[31:0];
          end
          ADDR_OUT_S30_DATA_0: begin
            rrdata <= int_out_s30[31:0];
          end
          ADDR_OUT_S31_DATA_0: begin
            rrdata <= int_out_s31[31:0];
          end
          ADDR_IN0_DATA_0: begin
            rrdata <= int_in0[31:0];
          end
          ADDR_IN0_DATA_1: begin
            rrdata <= int_in0[63:32];
          end
          ADDR_IN1_DATA_0: begin
            rrdata <= int_in1[31:0];
          end
          ADDR_IN1_DATA_1: begin
            rrdata <= int_in1[63:32];
          end
          ADDR_IN2_DATA_0: begin
            rrdata <= int_in2[31:0];
          end
          ADDR_IN2_DATA_1: begin
            rrdata <= int_in2[63:32];
          end
          ADDR_IN3_DATA_0: begin
            rrdata <= int_in3[31:0];
          end
          ADDR_IN3_DATA_1: begin
            rrdata <= int_in3[63:32];
          end
          ADDR_IN4_DATA_0: begin
            rrdata <= int_in4[31:0];
          end
          ADDR_IN4_DATA_1: begin
            rrdata <= int_in4[63:32];
          end
          ADDR_IN5_DATA_0: begin
            rrdata <= int_in5[31:0];
          end
          ADDR_IN5_DATA_1: begin
            rrdata <= int_in5[63:32];
          end
          ADDR_IN6_DATA_0: begin
            rrdata <= int_in6[31:0];
          end
          ADDR_IN6_DATA_1: begin
            rrdata <= int_in6[63:32];
          end
          ADDR_IN7_DATA_0: begin
            rrdata <= int_in7[31:0];
          end
          ADDR_IN7_DATA_1: begin
            rrdata <= int_in7[63:32];
          end
          ADDR_IN8_DATA_0: begin
            rrdata <= int_in8[31:0];
          end
          ADDR_IN8_DATA_1: begin
            rrdata <= int_in8[63:32];
          end
          ADDR_IN9_DATA_0: begin
            rrdata <= int_in9[31:0];
          end
          ADDR_IN9_DATA_1: begin
            rrdata <= int_in9[63:32];
          end
          ADDR_IN10_DATA_0: begin
            rrdata <= int_in10[31:0];
          end
          ADDR_IN10_DATA_1: begin
            rrdata <= int_in10[63:32];
          end
          ADDR_IN11_DATA_0: begin
            rrdata <= int_in11[31:0];
          end
          ADDR_IN11_DATA_1: begin
            rrdata <= int_in11[63:32];
          end
          ADDR_IN12_DATA_0: begin
            rrdata <= int_in12[31:0];
          end
          ADDR_IN12_DATA_1: begin
            rrdata <= int_in12[63:32];
          end
          ADDR_IN13_DATA_0: begin
            rrdata <= int_in13[31:0];
          end
          ADDR_IN13_DATA_1: begin
            rrdata <= int_in13[63:32];
          end
          ADDR_IN14_DATA_0: begin
            rrdata <= int_in14[31:0];
          end
          ADDR_IN14_DATA_1: begin
            rrdata <= int_in14[63:32];
          end
          ADDR_IN15_DATA_0: begin
            rrdata <= int_in15[31:0];
          end
          ADDR_IN15_DATA_1: begin
            rrdata <= int_in15[63:32];
          end
          ADDR_IN16_DATA_0: begin
            rrdata <= int_in16[31:0];
          end
          ADDR_IN16_DATA_1: begin
            rrdata <= int_in16[63:32];
          end
          ADDR_IN17_DATA_0: begin
            rrdata <= int_in17[31:0];
          end
          ADDR_IN17_DATA_1: begin
            rrdata <= int_in17[63:32];
          end
          ADDR_IN18_DATA_0: begin
            rrdata <= int_in18[31:0];
          end
          ADDR_IN18_DATA_1: begin
            rrdata <= int_in18[63:32];
          end
          ADDR_IN19_DATA_0: begin
            rrdata <= int_in19[31:0];
          end
          ADDR_IN19_DATA_1: begin
            rrdata <= int_in19[63:32];
          end
          ADDR_IN20_DATA_0: begin
            rrdata <= int_in20[31:0];
          end
          ADDR_IN20_DATA_1: begin
            rrdata <= int_in20[63:32];
          end
          ADDR_IN21_DATA_0: begin
            rrdata <= int_in21[31:0];
          end
          ADDR_IN21_DATA_1: begin
            rrdata <= int_in21[63:32];
          end
          ADDR_IN22_DATA_0: begin
            rrdata <= int_in22[31:0];
          end
          ADDR_IN22_DATA_1: begin
            rrdata <= int_in22[63:32];
          end
          ADDR_IN23_DATA_0: begin
            rrdata <= int_in23[31:0];
          end
          ADDR_IN23_DATA_1: begin
            rrdata <= int_in23[63:32];
          end
          ADDR_IN24_DATA_0: begin
            rrdata <= int_in24[31:0];
          end
          ADDR_IN24_DATA_1: begin
            rrdata <= int_in24[63:32];
          end
          ADDR_IN25_DATA_0: begin
            rrdata <= int_in25[31:0];
          end
          ADDR_IN25_DATA_1: begin
            rrdata <= int_in25[63:32];
          end
          ADDR_IN26_DATA_0: begin
            rrdata <= int_in26[31:0];
          end
          ADDR_IN26_DATA_1: begin
            rrdata <= int_in26[63:32];
          end
          ADDR_IN27_DATA_0: begin
            rrdata <= int_in27[31:0];
          end
          ADDR_IN27_DATA_1: begin
            rrdata <= int_in27[63:32];
          end
          ADDR_IN28_DATA_0: begin
            rrdata <= int_in28[31:0];
          end
          ADDR_IN28_DATA_1: begin
            rrdata <= int_in28[63:32];
          end
          ADDR_IN29_DATA_0: begin
            rrdata <= int_in29[31:0];
          end
          ADDR_IN29_DATA_1: begin
            rrdata <= int_in29[63:32];
          end
          ADDR_IN30_DATA_0: begin
            rrdata <= int_in30[31:0];
          end
          ADDR_IN30_DATA_1: begin
            rrdata <= int_in30[63:32];
          end
          ADDR_IN31_DATA_0: begin
            rrdata <= int_in31[31:0];
          end
          ADDR_IN31_DATA_1: begin
            rrdata <= int_in31[63:32];
          end
          ADDR_OUT0_DATA_0: begin
            rrdata <= int_out0[31:0];
          end
          ADDR_OUT0_DATA_1: begin
            rrdata <= int_out0[63:32];
          end
          ADDR_OUT1_DATA_0: begin
            rrdata <= int_out1[31:0];
          end
          ADDR_OUT1_DATA_1: begin
            rrdata <= int_out1[63:32];
          end
          ADDR_OUT2_DATA_0: begin
            rrdata <= int_out2[31:0];
          end
          ADDR_OUT2_DATA_1: begin
            rrdata <= int_out2[63:32];
          end
          ADDR_OUT3_DATA_0: begin
            rrdata <= int_out3[31:0];
          end
          ADDR_OUT3_DATA_1: begin
            rrdata <= int_out3[63:32];
          end
          ADDR_OUT4_DATA_0: begin
            rrdata <= int_out4[31:0];
          end
          ADDR_OUT4_DATA_1: begin
            rrdata <= int_out4[63:32];
          end
          ADDR_OUT5_DATA_0: begin
            rrdata <= int_out5[31:0];
          end
          ADDR_OUT5_DATA_1: begin
            rrdata <= int_out5[63:32];
          end
          ADDR_OUT6_DATA_0: begin
            rrdata <= int_out6[31:0];
          end
          ADDR_OUT6_DATA_1: begin
            rrdata <= int_out6[63:32];
          end
          ADDR_OUT7_DATA_0: begin
            rrdata <= int_out7[31:0];
          end
          ADDR_OUT7_DATA_1: begin
            rrdata <= int_out7[63:32];
          end
          ADDR_OUT8_DATA_0: begin
            rrdata <= int_out8[31:0];
          end
          ADDR_OUT8_DATA_1: begin
            rrdata <= int_out8[63:32];
          end
          ADDR_OUT9_DATA_0: begin
            rrdata <= int_out9[31:0];
          end
          ADDR_OUT9_DATA_1: begin
            rrdata <= int_out9[63:32];
          end
          ADDR_OUT10_DATA_0: begin
            rrdata <= int_out10[31:0];
          end
          ADDR_OUT10_DATA_1: begin
            rrdata <= int_out10[63:32];
          end
          ADDR_OUT11_DATA_0: begin
            rrdata <= int_out11[31:0];
          end
          ADDR_OUT11_DATA_1: begin
            rrdata <= int_out11[63:32];
          end
          ADDR_OUT12_DATA_0: begin
            rrdata <= int_out12[31:0];
          end
          ADDR_OUT12_DATA_1: begin
            rrdata <= int_out12[63:32];
          end
          ADDR_OUT13_DATA_0: begin
            rrdata <= int_out13[31:0];
          end
          ADDR_OUT13_DATA_1: begin
            rrdata <= int_out13[63:32];
          end
          ADDR_OUT14_DATA_0: begin
            rrdata <= int_out14[31:0];
          end
          ADDR_OUT14_DATA_1: begin
            rrdata <= int_out14[63:32];
          end
          ADDR_OUT15_DATA_0: begin
            rrdata <= int_out15[31:0];
          end
          ADDR_OUT15_DATA_1: begin
            rrdata <= int_out15[63:32];
          end
          ADDR_OUT16_DATA_0: begin
            rrdata <= int_out16[31:0];
          end
          ADDR_OUT16_DATA_1: begin
            rrdata <= int_out16[63:32];
          end
          ADDR_OUT17_DATA_0: begin
            rrdata <= int_out17[31:0];
          end
          ADDR_OUT17_DATA_1: begin
            rrdata <= int_out17[63:32];
          end
          ADDR_OUT18_DATA_0: begin
            rrdata <= int_out18[31:0];
          end
          ADDR_OUT18_DATA_1: begin
            rrdata <= int_out18[63:32];
          end
          ADDR_OUT19_DATA_0: begin
            rrdata <= int_out19[31:0];
          end
          ADDR_OUT19_DATA_1: begin
            rrdata <= int_out19[63:32];
          end
          ADDR_OUT20_DATA_0: begin
            rrdata <= int_out20[31:0];
          end
          ADDR_OUT20_DATA_1: begin
            rrdata <= int_out20[63:32];
          end
          ADDR_OUT21_DATA_0: begin
            rrdata <= int_out21[31:0];
          end
          ADDR_OUT21_DATA_1: begin
            rrdata <= int_out21[63:32];
          end
          ADDR_OUT22_DATA_0: begin
            rrdata <= int_out22[31:0];
          end
          ADDR_OUT22_DATA_1: begin
            rrdata <= int_out22[63:32];
          end
          ADDR_OUT23_DATA_0: begin
            rrdata <= int_out23[31:0];
          end
          ADDR_OUT23_DATA_1: begin
            rrdata <= int_out23[63:32];
          end
          ADDR_OUT24_DATA_0: begin
            rrdata <= int_out24[31:0];
          end
          ADDR_OUT24_DATA_1: begin
            rrdata <= int_out24[63:32];
          end
          ADDR_OUT25_DATA_0: begin
            rrdata <= int_out25[31:0];
          end
          ADDR_OUT25_DATA_1: begin
            rrdata <= int_out25[63:32];
          end
          ADDR_OUT26_DATA_0: begin
            rrdata <= int_out26[31:0];
          end
          ADDR_OUT26_DATA_1: begin
            rrdata <= int_out26[63:32];
          end
          ADDR_OUT27_DATA_0: begin
            rrdata <= int_out27[31:0];
          end
          ADDR_OUT27_DATA_1: begin
            rrdata <= int_out27[63:32];
          end
          ADDR_OUT28_DATA_0: begin
            rrdata <= int_out28[31:0];
          end
          ADDR_OUT28_DATA_1: begin
            rrdata <= int_out28[63:32];
          end
          ADDR_OUT29_DATA_0: begin
            rrdata <= int_out29[31:0];
          end
          ADDR_OUT29_DATA_1: begin
            rrdata <= int_out29[63:32];
          end
          ADDR_OUT30_DATA_0: begin
            rrdata <= int_out30[31:0];
          end
          ADDR_OUT30_DATA_1: begin
            rrdata <= int_out30[63:32];
          end
          ADDR_OUT31_DATA_0: begin
            rrdata <= int_out31[31:0];
          end
          ADDR_OUT31_DATA_1: begin
            rrdata <= int_out31[63:32];
          end
        endcase
      end 
    end 
  end

  assign interrupt = int_gie & |int_isr;
  assign ap_start = int_ap_start;
  assign in_s0 = int_in_s0;
  assign in_s1 = int_in_s1;
  assign in_s2 = int_in_s2;
  assign in_s3 = int_in_s3;
  assign in_s4 = int_in_s4;
  assign in_s5 = int_in_s5;
  assign in_s6 = int_in_s6;
  assign in_s7 = int_in_s7;
  assign in_s8 = int_in_s8;
  assign in_s9 = int_in_s9;
  assign in_s10 = int_in_s10;
  assign in_s11 = int_in_s11;
  assign in_s12 = int_in_s12;
  assign in_s13 = int_in_s13;
  assign in_s14 = int_in_s14;
  assign in_s15 = int_in_s15;
  assign in_s16 = int_in_s16;
  assign in_s17 = int_in_s17;
  assign in_s18 = int_in_s18;
  assign in_s19 = int_in_s19;
  assign in_s20 = int_in_s20;
  assign in_s21 = int_in_s21;
  assign in_s22 = int_in_s22;
  assign in_s23 = int_in_s23;
  assign in_s24 = int_in_s24;
  assign in_s25 = int_in_s25;
  assign in_s26 = int_in_s26;
  assign in_s27 = int_in_s27;
  assign in_s28 = int_in_s28;
  assign in_s29 = int_in_s29;
  assign in_s30 = int_in_s30;
  assign in_s31 = int_in_s31;
  assign out_s0 = int_out_s0;
  assign out_s1 = int_out_s1;
  assign out_s2 = int_out_s2;
  assign out_s3 = int_out_s3;
  assign out_s4 = int_out_s4;
  assign out_s5 = int_out_s5;
  assign out_s6 = int_out_s6;
  assign out_s7 = int_out_s7;
  assign out_s8 = int_out_s8;
  assign out_s9 = int_out_s9;
  assign out_s10 = int_out_s10;
  assign out_s11 = int_out_s11;
  assign out_s12 = int_out_s12;
  assign out_s13 = int_out_s13;
  assign out_s14 = int_out_s14;
  assign out_s15 = int_out_s15;
  assign out_s16 = int_out_s16;
  assign out_s17 = int_out_s17;
  assign out_s18 = int_out_s18;
  assign out_s19 = int_out_s19;
  assign out_s20 = int_out_s20;
  assign out_s21 = int_out_s21;
  assign out_s22 = int_out_s22;
  assign out_s23 = int_out_s23;
  assign out_s24 = int_out_s24;
  assign out_s25 = int_out_s25;
  assign out_s26 = int_out_s26;
  assign out_s27 = int_out_s27;
  assign out_s28 = int_out_s28;
  assign out_s29 = int_out_s29;
  assign out_s30 = int_out_s30;
  assign out_s31 = int_out_s31;
  assign in0 = int_in0;
  assign out0 = int_out0;
  assign in1 = int_in1;
  assign out1 = int_out1;
  assign in2 = int_in2;
  assign out2 = int_out2;
  assign in3 = int_in3;
  assign out3 = int_out3;
  assign in4 = int_in4;
  assign out4 = int_out4;
  assign in5 = int_in5;
  assign out5 = int_out5;
  assign in6 = int_in6;
  assign out6 = int_out6;
  assign in7 = int_in7;
  assign out7 = int_out7;
  assign in8 = int_in8;
  assign out8 = int_out8;
  assign in9 = int_in9;
  assign out9 = int_out9;
  assign in10 = int_in10;
  assign out10 = int_out10;
  assign in11 = int_in11;
  assign out11 = int_out11;
  assign in12 = int_in12;
  assign out12 = int_out12;
  assign in13 = int_in13;
  assign out13 = int_out13;
  assign in14 = int_in14;
  assign out14 = int_out14;
  assign in15 = int_in15;
  assign out15 = int_out15;
  assign in16 = int_in16;
  assign out16 = int_out16;
  assign in17 = int_in17;
  assign out17 = int_out17;
  assign in18 = int_in18;
  assign out18 = int_out18;
  assign in19 = int_in19;
  assign out19 = int_out19;
  assign in20 = int_in20;
  assign out20 = int_out20;
  assign in21 = int_in21;
  assign out21 = int_out21;
  assign in22 = int_in22;
  assign out22 = int_out22;
  assign in23 = int_in23;
  assign out23 = int_out23;
  assign in24 = int_in24;
  assign out24 = int_out24;
  assign in25 = int_in25;
  assign out25 = int_out25;
  assign in26 = int_in26;
  assign out26 = int_out26;
  assign in27 = int_in27;
  assign out27 = int_out27;
  assign in28 = int_in28;
  assign out28 = int_out28;
  assign in29 = int_in29;
  assign out29 = int_out29;
  assign in30 = int_in30;
  assign out30 = int_out30;
  assign in31 = int_in31;
  assign out31 = int_out31;

  always @(posedge aclk) begin
    if(areset) begin
      int_ap_start <= 1'b0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_AP_CTRL) && wstrb[0] && wdata[0]) begin
          int_ap_start <= 1'b1;
        end else if(ap_ready) begin
          int_ap_start <= int_auto_restart;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_ap_done <= 1'b0;
    end else begin
      if(aclk_en) begin
        if(ap_done) begin
          int_ap_done <= 1'b1;
        end else if(ar_hs && (raddr == ADDR_AP_CTRL)) begin
          int_ap_done <= 1'b0;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_ap_idle <= 1'b1;
    end else begin
      if(aclk_en) begin
        int_ap_idle <= ap_idle;
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_ap_ready <= 1'b0;
    end else begin
      if(aclk_en) begin
        int_ap_ready <= ap_ready;
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_auto_restart <= 1'b0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_AP_CTRL) && wstrb[0]) begin
          int_auto_restart <= wdata[7];
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_gie <= 1'b0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_GIE) && wstrb[0]) begin
          int_gie <= wdata[0];
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_ier <= 2'b0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IER) && wstrb[0]) begin
          int_ier <= wdata[1:0];
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_isr[0] <= 1'b0;
    end else begin
      if(aclk_en) begin
        if(int_ier[0] & ap_done) begin
          int_isr[0] <= 1'b1;
        end else if(w_hs && (waddr == ADDR_ISR) && wstrb[0]) begin
          int_isr[0] <= int_isr[0] ^ wdata[0];
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_isr[1] <= 1'b0;
    end else begin
      if(aclk_en) begin
        if(int_ier[1] & ap_ready) begin
          int_isr[1] <= 1'b1;
        end else if(w_hs && (waddr == ADDR_ISR) && wstrb[0]) begin
          int_isr[1] <= int_isr[1] ^ wdata[1];
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s0[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S0_DATA_0)) begin
          int_in_s0[31:0] <= wdata[31:0] & wmask | int_in_s0[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s1[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S1_DATA_0)) begin
          int_in_s1[31:0] <= wdata[31:0] & wmask | int_in_s1[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s2[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S2_DATA_0)) begin
          int_in_s2[31:0] <= wdata[31:0] & wmask | int_in_s2[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s3[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S3_DATA_0)) begin
          int_in_s3[31:0] <= wdata[31:0] & wmask | int_in_s3[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s4[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S4_DATA_0)) begin
          int_in_s4[31:0] <= wdata[31:0] & wmask | int_in_s4[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s5[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S5_DATA_0)) begin
          int_in_s5[31:0] <= wdata[31:0] & wmask | int_in_s5[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s6[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S6_DATA_0)) begin
          int_in_s6[31:0] <= wdata[31:0] & wmask | int_in_s6[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s7[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S7_DATA_0)) begin
          int_in_s7[31:0] <= wdata[31:0] & wmask | int_in_s7[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s8[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S8_DATA_0)) begin
          int_in_s8[31:0] <= wdata[31:0] & wmask | int_in_s8[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s9[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S9_DATA_0)) begin
          int_in_s9[31:0] <= wdata[31:0] & wmask | int_in_s9[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s10[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S10_DATA_0)) begin
          int_in_s10[31:0] <= wdata[31:0] & wmask | int_in_s10[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s11[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S11_DATA_0)) begin
          int_in_s11[31:0] <= wdata[31:0] & wmask | int_in_s11[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s12[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S12_DATA_0)) begin
          int_in_s12[31:0] <= wdata[31:0] & wmask | int_in_s12[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s13[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S13_DATA_0)) begin
          int_in_s13[31:0] <= wdata[31:0] & wmask | int_in_s13[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s14[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S14_DATA_0)) begin
          int_in_s14[31:0] <= wdata[31:0] & wmask | int_in_s14[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s15[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S15_DATA_0)) begin
          int_in_s15[31:0] <= wdata[31:0] & wmask | int_in_s15[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s16[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S16_DATA_0)) begin
          int_in_s16[31:0] <= wdata[31:0] & wmask | int_in_s16[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s17[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S17_DATA_0)) begin
          int_in_s17[31:0] <= wdata[31:0] & wmask | int_in_s17[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s18[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S18_DATA_0)) begin
          int_in_s18[31:0] <= wdata[31:0] & wmask | int_in_s18[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s19[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S19_DATA_0)) begin
          int_in_s19[31:0] <= wdata[31:0] & wmask | int_in_s19[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s20[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S20_DATA_0)) begin
          int_in_s20[31:0] <= wdata[31:0] & wmask | int_in_s20[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s21[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S21_DATA_0)) begin
          int_in_s21[31:0] <= wdata[31:0] & wmask | int_in_s21[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s22[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S22_DATA_0)) begin
          int_in_s22[31:0] <= wdata[31:0] & wmask | int_in_s22[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s23[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S23_DATA_0)) begin
          int_in_s23[31:0] <= wdata[31:0] & wmask | int_in_s23[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s24[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S24_DATA_0)) begin
          int_in_s24[31:0] <= wdata[31:0] & wmask | int_in_s24[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s25[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S25_DATA_0)) begin
          int_in_s25[31:0] <= wdata[31:0] & wmask | int_in_s25[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s26[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S26_DATA_0)) begin
          int_in_s26[31:0] <= wdata[31:0] & wmask | int_in_s26[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s27[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S27_DATA_0)) begin
          int_in_s27[31:0] <= wdata[31:0] & wmask | int_in_s27[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s28[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S28_DATA_0)) begin
          int_in_s28[31:0] <= wdata[31:0] & wmask | int_in_s28[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s29[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S29_DATA_0)) begin
          int_in_s29[31:0] <= wdata[31:0] & wmask | int_in_s29[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s30[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S30_DATA_0)) begin
          int_in_s30[31:0] <= wdata[31:0] & wmask | int_in_s30[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in_s31[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN_S31_DATA_0)) begin
          int_in_s31[31:0] <= wdata[31:0] & wmask | int_in_s31[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s0[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S0_DATA_0)) begin
          int_out_s0[31:0] <= wdata[31:0] & wmask | int_out_s0[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s1[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S1_DATA_0)) begin
          int_out_s1[31:0] <= wdata[31:0] & wmask | int_out_s1[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s2[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S2_DATA_0)) begin
          int_out_s2[31:0] <= wdata[31:0] & wmask | int_out_s2[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s3[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S3_DATA_0)) begin
          int_out_s3[31:0] <= wdata[31:0] & wmask | int_out_s3[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s4[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S4_DATA_0)) begin
          int_out_s4[31:0] <= wdata[31:0] & wmask | int_out_s4[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s5[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S5_DATA_0)) begin
          int_out_s5[31:0] <= wdata[31:0] & wmask | int_out_s5[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s6[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S6_DATA_0)) begin
          int_out_s6[31:0] <= wdata[31:0] & wmask | int_out_s6[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s7[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S7_DATA_0)) begin
          int_out_s7[31:0] <= wdata[31:0] & wmask | int_out_s7[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s8[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S8_DATA_0)) begin
          int_out_s8[31:0] <= wdata[31:0] & wmask | int_out_s8[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s9[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S9_DATA_0)) begin
          int_out_s9[31:0] <= wdata[31:0] & wmask | int_out_s9[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s10[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S10_DATA_0)) begin
          int_out_s10[31:0] <= wdata[31:0] & wmask | int_out_s10[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s11[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S11_DATA_0)) begin
          int_out_s11[31:0] <= wdata[31:0] & wmask | int_out_s11[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s12[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S12_DATA_0)) begin
          int_out_s12[31:0] <= wdata[31:0] & wmask | int_out_s12[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s13[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S13_DATA_0)) begin
          int_out_s13[31:0] <= wdata[31:0] & wmask | int_out_s13[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s14[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S14_DATA_0)) begin
          int_out_s14[31:0] <= wdata[31:0] & wmask | int_out_s14[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s15[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S15_DATA_0)) begin
          int_out_s15[31:0] <= wdata[31:0] & wmask | int_out_s15[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s16[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S16_DATA_0)) begin
          int_out_s16[31:0] <= wdata[31:0] & wmask | int_out_s16[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s17[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S17_DATA_0)) begin
          int_out_s17[31:0] <= wdata[31:0] & wmask | int_out_s17[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s18[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S18_DATA_0)) begin
          int_out_s18[31:0] <= wdata[31:0] & wmask | int_out_s18[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s19[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S19_DATA_0)) begin
          int_out_s19[31:0] <= wdata[31:0] & wmask | int_out_s19[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s20[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S20_DATA_0)) begin
          int_out_s20[31:0] <= wdata[31:0] & wmask | int_out_s20[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s21[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S21_DATA_0)) begin
          int_out_s21[31:0] <= wdata[31:0] & wmask | int_out_s21[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s22[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S22_DATA_0)) begin
          int_out_s22[31:0] <= wdata[31:0] & wmask | int_out_s22[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s23[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S23_DATA_0)) begin
          int_out_s23[31:0] <= wdata[31:0] & wmask | int_out_s23[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s24[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S24_DATA_0)) begin
          int_out_s24[31:0] <= wdata[31:0] & wmask | int_out_s24[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s25[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S25_DATA_0)) begin
          int_out_s25[31:0] <= wdata[31:0] & wmask | int_out_s25[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s26[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S26_DATA_0)) begin
          int_out_s26[31:0] <= wdata[31:0] & wmask | int_out_s26[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s27[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S27_DATA_0)) begin
          int_out_s27[31:0] <= wdata[31:0] & wmask | int_out_s27[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s28[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S28_DATA_0)) begin
          int_out_s28[31:0] <= wdata[31:0] & wmask | int_out_s28[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s29[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S29_DATA_0)) begin
          int_out_s29[31:0] <= wdata[31:0] & wmask | int_out_s29[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s30[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S30_DATA_0)) begin
          int_out_s30[31:0] <= wdata[31:0] & wmask | int_out_s30[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out_s31[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT_S31_DATA_0)) begin
          int_out_s31[31:0] <= wdata[31:0] & wmask | int_out_s31[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in0[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN0_DATA_0)) begin
          int_in0[31:0] <= wdata[31:0] & wmask | int_in0[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in0[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN0_DATA_1)) begin
          int_in0[63:32] <= wdata[31:0] & wmask | int_in0[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out0[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT0_DATA_0)) begin
          int_out0[31:0] <= wdata[31:0] & wmask | int_out0[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out0[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT0_DATA_1)) begin
          int_out0[63:32] <= wdata[31:0] & wmask | int_out0[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in1[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN1_DATA_0)) begin
          int_in1[31:0] <= wdata[31:0] & wmask | int_in1[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in1[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN1_DATA_1)) begin
          int_in1[63:32] <= wdata[31:0] & wmask | int_in1[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out1[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT1_DATA_0)) begin
          int_out1[31:0] <= wdata[31:0] & wmask | int_out1[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out1[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT1_DATA_1)) begin
          int_out1[63:32] <= wdata[31:0] & wmask | int_out1[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in2[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN2_DATA_0)) begin
          int_in2[31:0] <= wdata[31:0] & wmask | int_in2[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in2[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN2_DATA_1)) begin
          int_in2[63:32] <= wdata[31:0] & wmask | int_in2[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out2[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT2_DATA_0)) begin
          int_out2[31:0] <= wdata[31:0] & wmask | int_out2[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out2[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT2_DATA_1)) begin
          int_out2[63:32] <= wdata[31:0] & wmask | int_out2[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in3[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN3_DATA_0)) begin
          int_in3[31:0] <= wdata[31:0] & wmask | int_in3[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in3[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN3_DATA_1)) begin
          int_in3[63:32] <= wdata[31:0] & wmask | int_in3[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out3[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT3_DATA_0)) begin
          int_out3[31:0] <= wdata[31:0] & wmask | int_out3[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out3[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT3_DATA_1)) begin
          int_out3[63:32] <= wdata[31:0] & wmask | int_out3[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in4[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN4_DATA_0)) begin
          int_in4[31:0] <= wdata[31:0] & wmask | int_in4[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in4[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN4_DATA_1)) begin
          int_in4[63:32] <= wdata[31:0] & wmask | int_in4[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out4[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT4_DATA_0)) begin
          int_out4[31:0] <= wdata[31:0] & wmask | int_out4[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out4[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT4_DATA_1)) begin
          int_out4[63:32] <= wdata[31:0] & wmask | int_out4[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in5[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN5_DATA_0)) begin
          int_in5[31:0] <= wdata[31:0] & wmask | int_in5[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in5[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN5_DATA_1)) begin
          int_in5[63:32] <= wdata[31:0] & wmask | int_in5[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out5[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT5_DATA_0)) begin
          int_out5[31:0] <= wdata[31:0] & wmask | int_out5[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out5[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT5_DATA_1)) begin
          int_out5[63:32] <= wdata[31:0] & wmask | int_out5[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in6[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN6_DATA_0)) begin
          int_in6[31:0] <= wdata[31:0] & wmask | int_in6[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in6[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN6_DATA_1)) begin
          int_in6[63:32] <= wdata[31:0] & wmask | int_in6[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out6[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT6_DATA_0)) begin
          int_out6[31:0] <= wdata[31:0] & wmask | int_out6[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out6[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT6_DATA_1)) begin
          int_out6[63:32] <= wdata[31:0] & wmask | int_out6[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in7[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN7_DATA_0)) begin
          int_in7[31:0] <= wdata[31:0] & wmask | int_in7[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in7[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN7_DATA_1)) begin
          int_in7[63:32] <= wdata[31:0] & wmask | int_in7[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out7[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT7_DATA_0)) begin
          int_out7[31:0] <= wdata[31:0] & wmask | int_out7[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out7[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT7_DATA_1)) begin
          int_out7[63:32] <= wdata[31:0] & wmask | int_out7[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in8[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN8_DATA_0)) begin
          int_in8[31:0] <= wdata[31:0] & wmask | int_in8[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in8[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN8_DATA_1)) begin
          int_in8[63:32] <= wdata[31:0] & wmask | int_in8[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out8[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT8_DATA_0)) begin
          int_out8[31:0] <= wdata[31:0] & wmask | int_out8[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out8[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT8_DATA_1)) begin
          int_out8[63:32] <= wdata[31:0] & wmask | int_out8[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in9[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN9_DATA_0)) begin
          int_in9[31:0] <= wdata[31:0] & wmask | int_in9[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in9[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN9_DATA_1)) begin
          int_in9[63:32] <= wdata[31:0] & wmask | int_in9[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out9[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT9_DATA_0)) begin
          int_out9[31:0] <= wdata[31:0] & wmask | int_out9[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out9[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT9_DATA_1)) begin
          int_out9[63:32] <= wdata[31:0] & wmask | int_out9[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in10[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN10_DATA_0)) begin
          int_in10[31:0] <= wdata[31:0] & wmask | int_in10[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in10[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN10_DATA_1)) begin
          int_in10[63:32] <= wdata[31:0] & wmask | int_in10[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out10[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT10_DATA_0)) begin
          int_out10[31:0] <= wdata[31:0] & wmask | int_out10[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out10[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT10_DATA_1)) begin
          int_out10[63:32] <= wdata[31:0] & wmask | int_out10[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in11[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN11_DATA_0)) begin
          int_in11[31:0] <= wdata[31:0] & wmask | int_in11[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in11[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN11_DATA_1)) begin
          int_in11[63:32] <= wdata[31:0] & wmask | int_in11[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out11[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT11_DATA_0)) begin
          int_out11[31:0] <= wdata[31:0] & wmask | int_out11[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out11[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT11_DATA_1)) begin
          int_out11[63:32] <= wdata[31:0] & wmask | int_out11[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in12[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN12_DATA_0)) begin
          int_in12[31:0] <= wdata[31:0] & wmask | int_in12[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in12[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN12_DATA_1)) begin
          int_in12[63:32] <= wdata[31:0] & wmask | int_in12[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out12[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT12_DATA_0)) begin
          int_out12[31:0] <= wdata[31:0] & wmask | int_out12[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out12[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT12_DATA_1)) begin
          int_out12[63:32] <= wdata[31:0] & wmask | int_out12[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in13[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN13_DATA_0)) begin
          int_in13[31:0] <= wdata[31:0] & wmask | int_in13[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in13[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN13_DATA_1)) begin
          int_in13[63:32] <= wdata[31:0] & wmask | int_in13[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out13[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT13_DATA_0)) begin
          int_out13[31:0] <= wdata[31:0] & wmask | int_out13[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out13[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT13_DATA_1)) begin
          int_out13[63:32] <= wdata[31:0] & wmask | int_out13[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in14[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN14_DATA_0)) begin
          int_in14[31:0] <= wdata[31:0] & wmask | int_in14[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in14[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN14_DATA_1)) begin
          int_in14[63:32] <= wdata[31:0] & wmask | int_in14[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out14[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT14_DATA_0)) begin
          int_out14[31:0] <= wdata[31:0] & wmask | int_out14[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out14[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT14_DATA_1)) begin
          int_out14[63:32] <= wdata[31:0] & wmask | int_out14[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in15[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN15_DATA_0)) begin
          int_in15[31:0] <= wdata[31:0] & wmask | int_in15[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in15[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN15_DATA_1)) begin
          int_in15[63:32] <= wdata[31:0] & wmask | int_in15[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out15[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT15_DATA_0)) begin
          int_out15[31:0] <= wdata[31:0] & wmask | int_out15[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out15[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT15_DATA_1)) begin
          int_out15[63:32] <= wdata[31:0] & wmask | int_out15[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in16[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN16_DATA_0)) begin
          int_in16[31:0] <= wdata[31:0] & wmask | int_in16[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in16[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN16_DATA_1)) begin
          int_in16[63:32] <= wdata[31:0] & wmask | int_in16[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out16[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT16_DATA_0)) begin
          int_out16[31:0] <= wdata[31:0] & wmask | int_out16[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out16[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT16_DATA_1)) begin
          int_out16[63:32] <= wdata[31:0] & wmask | int_out16[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in17[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN17_DATA_0)) begin
          int_in17[31:0] <= wdata[31:0] & wmask | int_in17[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in17[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN17_DATA_1)) begin
          int_in17[63:32] <= wdata[31:0] & wmask | int_in17[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out17[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT17_DATA_0)) begin
          int_out17[31:0] <= wdata[31:0] & wmask | int_out17[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out17[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT17_DATA_1)) begin
          int_out17[63:32] <= wdata[31:0] & wmask | int_out17[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in18[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN18_DATA_0)) begin
          int_in18[31:0] <= wdata[31:0] & wmask | int_in18[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in18[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN18_DATA_1)) begin
          int_in18[63:32] <= wdata[31:0] & wmask | int_in18[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out18[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT18_DATA_0)) begin
          int_out18[31:0] <= wdata[31:0] & wmask | int_out18[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out18[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT18_DATA_1)) begin
          int_out18[63:32] <= wdata[31:0] & wmask | int_out18[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in19[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN19_DATA_0)) begin
          int_in19[31:0] <= wdata[31:0] & wmask | int_in19[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in19[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN19_DATA_1)) begin
          int_in19[63:32] <= wdata[31:0] & wmask | int_in19[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out19[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT19_DATA_0)) begin
          int_out19[31:0] <= wdata[31:0] & wmask | int_out19[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out19[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT19_DATA_1)) begin
          int_out19[63:32] <= wdata[31:0] & wmask | int_out19[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in20[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN20_DATA_0)) begin
          int_in20[31:0] <= wdata[31:0] & wmask | int_in20[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in20[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN20_DATA_1)) begin
          int_in20[63:32] <= wdata[31:0] & wmask | int_in20[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out20[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT20_DATA_0)) begin
          int_out20[31:0] <= wdata[31:0] & wmask | int_out20[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out20[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT20_DATA_1)) begin
          int_out20[63:32] <= wdata[31:0] & wmask | int_out20[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in21[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN21_DATA_0)) begin
          int_in21[31:0] <= wdata[31:0] & wmask | int_in21[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in21[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN21_DATA_1)) begin
          int_in21[63:32] <= wdata[31:0] & wmask | int_in21[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out21[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT21_DATA_0)) begin
          int_out21[31:0] <= wdata[31:0] & wmask | int_out21[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out21[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT21_DATA_1)) begin
          int_out21[63:32] <= wdata[31:0] & wmask | int_out21[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in22[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN22_DATA_0)) begin
          int_in22[31:0] <= wdata[31:0] & wmask | int_in22[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in22[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN22_DATA_1)) begin
          int_in22[63:32] <= wdata[31:0] & wmask | int_in22[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out22[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT22_DATA_0)) begin
          int_out22[31:0] <= wdata[31:0] & wmask | int_out22[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out22[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT22_DATA_1)) begin
          int_out22[63:32] <= wdata[31:0] & wmask | int_out22[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in23[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN23_DATA_0)) begin
          int_in23[31:0] <= wdata[31:0] & wmask | int_in23[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in23[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN23_DATA_1)) begin
          int_in23[63:32] <= wdata[31:0] & wmask | int_in23[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out23[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT23_DATA_0)) begin
          int_out23[31:0] <= wdata[31:0] & wmask | int_out23[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out23[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT23_DATA_1)) begin
          int_out23[63:32] <= wdata[31:0] & wmask | int_out23[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in24[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN24_DATA_0)) begin
          int_in24[31:0] <= wdata[31:0] & wmask | int_in24[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in24[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN24_DATA_1)) begin
          int_in24[63:32] <= wdata[31:0] & wmask | int_in24[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out24[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT24_DATA_0)) begin
          int_out24[31:0] <= wdata[31:0] & wmask | int_out24[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out24[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT24_DATA_1)) begin
          int_out24[63:32] <= wdata[31:0] & wmask | int_out24[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in25[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN25_DATA_0)) begin
          int_in25[31:0] <= wdata[31:0] & wmask | int_in25[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in25[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN25_DATA_1)) begin
          int_in25[63:32] <= wdata[31:0] & wmask | int_in25[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out25[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT25_DATA_0)) begin
          int_out25[31:0] <= wdata[31:0] & wmask | int_out25[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out25[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT25_DATA_1)) begin
          int_out25[63:32] <= wdata[31:0] & wmask | int_out25[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in26[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN26_DATA_0)) begin
          int_in26[31:0] <= wdata[31:0] & wmask | int_in26[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in26[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN26_DATA_1)) begin
          int_in26[63:32] <= wdata[31:0] & wmask | int_in26[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out26[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT26_DATA_0)) begin
          int_out26[31:0] <= wdata[31:0] & wmask | int_out26[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out26[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT26_DATA_1)) begin
          int_out26[63:32] <= wdata[31:0] & wmask | int_out26[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in27[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN27_DATA_0)) begin
          int_in27[31:0] <= wdata[31:0] & wmask | int_in27[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in27[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN27_DATA_1)) begin
          int_in27[63:32] <= wdata[31:0] & wmask | int_in27[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out27[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT27_DATA_0)) begin
          int_out27[31:0] <= wdata[31:0] & wmask | int_out27[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out27[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT27_DATA_1)) begin
          int_out27[63:32] <= wdata[31:0] & wmask | int_out27[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in28[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN28_DATA_0)) begin
          int_in28[31:0] <= wdata[31:0] & wmask | int_in28[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in28[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN28_DATA_1)) begin
          int_in28[63:32] <= wdata[31:0] & wmask | int_in28[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out28[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT28_DATA_0)) begin
          int_out28[31:0] <= wdata[31:0] & wmask | int_out28[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out28[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT28_DATA_1)) begin
          int_out28[63:32] <= wdata[31:0] & wmask | int_out28[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in29[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN29_DATA_0)) begin
          int_in29[31:0] <= wdata[31:0] & wmask | int_in29[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in29[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN29_DATA_1)) begin
          int_in29[63:32] <= wdata[31:0] & wmask | int_in29[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out29[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT29_DATA_0)) begin
          int_out29[31:0] <= wdata[31:0] & wmask | int_out29[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out29[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT29_DATA_1)) begin
          int_out29[63:32] <= wdata[31:0] & wmask | int_out29[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in30[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN30_DATA_0)) begin
          int_in30[31:0] <= wdata[31:0] & wmask | int_in30[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in30[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN30_DATA_1)) begin
          int_in30[63:32] <= wdata[31:0] & wmask | int_in30[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out30[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT30_DATA_0)) begin
          int_out30[31:0] <= wdata[31:0] & wmask | int_out30[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out30[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT30_DATA_1)) begin
          int_out30[63:32] <= wdata[31:0] & wmask | int_out30[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in31[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN31_DATA_0)) begin
          int_in31[31:0] <= wdata[31:0] & wmask | int_in31[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_in31[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_IN31_DATA_1)) begin
          int_in31[63:32] <= wdata[31:0] & wmask | int_in31[63:32] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out31[31:0] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT31_DATA_0)) begin
          int_out31[31:0] <= wdata[31:0] & wmask | int_out31[31:0] & ~wmask;
        end 
      end 
    end
  end


  always @(posedge aclk) begin
    if(areset) begin
      int_out31[63:32] <= 32'd0;
    end else begin
      if(aclk_en) begin
        if(w_hs && (waddr == ADDR_OUT31_DATA_1)) begin
          int_out31[63:32] <= wdata[31:0] & wmask | int_out31[63:32] & ~wmask;
        end 
      end 
    end
  end


  initial begin
    wstate = WRRESET;
    wnext = 0;
    waddr = 0;
    rstate = RDRESET;
    rnext = 0;
    rrdata = 0;
    int_ap_idle = 1'b1;
    int_ap_ready = 0;
    int_ap_done = 0;
    int_ap_start = 0;
    int_auto_restart = 0;
    int_gie = 0;
    int_ier = 0;
    int_isr = 0;
    int_in_s0 = 0;
    int_in_s1 = 0;
    int_in_s2 = 0;
    int_in_s3 = 0;
    int_in_s4 = 0;
    int_in_s5 = 0;
    int_in_s6 = 0;
    int_in_s7 = 0;
    int_in_s8 = 0;
    int_in_s9 = 0;
    int_in_s10 = 0;
    int_in_s11 = 0;
    int_in_s12 = 0;
    int_in_s13 = 0;
    int_in_s14 = 0;
    int_in_s15 = 0;
    int_in_s16 = 0;
    int_in_s17 = 0;
    int_in_s18 = 0;
    int_in_s19 = 0;
    int_in_s20 = 0;
    int_in_s21 = 0;
    int_in_s22 = 0;
    int_in_s23 = 0;
    int_in_s24 = 0;
    int_in_s25 = 0;
    int_in_s26 = 0;
    int_in_s27 = 0;
    int_in_s28 = 0;
    int_in_s29 = 0;
    int_in_s30 = 0;
    int_in_s31 = 0;
    int_out_s0 = 0;
    int_out_s1 = 0;
    int_out_s2 = 0;
    int_out_s3 = 0;
    int_out_s4 = 0;
    int_out_s5 = 0;
    int_out_s6 = 0;
    int_out_s7 = 0;
    int_out_s8 = 0;
    int_out_s9 = 0;
    int_out_s10 = 0;
    int_out_s11 = 0;
    int_out_s12 = 0;
    int_out_s13 = 0;
    int_out_s14 = 0;
    int_out_s15 = 0;
    int_out_s16 = 0;
    int_out_s17 = 0;
    int_out_s18 = 0;
    int_out_s19 = 0;
    int_out_s20 = 0;
    int_out_s21 = 0;
    int_out_s22 = 0;
    int_out_s23 = 0;
    int_out_s24 = 0;
    int_out_s25 = 0;
    int_out_s26 = 0;
    int_out_s27 = 0;
    int_out_s28 = 0;
    int_out_s29 = 0;
    int_out_s30 = 0;
    int_out_s31 = 0;
    int_in0 = 0;
    int_out0 = 0;
    int_in1 = 0;
    int_out1 = 0;
    int_in2 = 0;
    int_out2 = 0;
    int_in3 = 0;
    int_out3 = 0;
    int_in4 = 0;
    int_out4 = 0;
    int_in5 = 0;
    int_out5 = 0;
    int_in6 = 0;
    int_out6 = 0;
    int_in7 = 0;
    int_out7 = 0;
    int_in8 = 0;
    int_out8 = 0;
    int_in9 = 0;
    int_out9 = 0;
    int_in10 = 0;
    int_out10 = 0;
    int_in11 = 0;
    int_out11 = 0;
    int_in12 = 0;
    int_out12 = 0;
    int_in13 = 0;
    int_out13 = 0;
    int_in14 = 0;
    int_out14 = 0;
    int_in15 = 0;
    int_out15 = 0;
    int_in16 = 0;
    int_out16 = 0;
    int_in17 = 0;
    int_out17 = 0;
    int_in18 = 0;
    int_out18 = 0;
    int_in19 = 0;
    int_out19 = 0;
    int_in20 = 0;
    int_out20 = 0;
    int_in21 = 0;
    int_out21 = 0;
    int_in22 = 0;
    int_out22 = 0;
    int_in23 = 0;
    int_out23 = 0;
    int_in24 = 0;
    int_out24 = 0;
    int_in25 = 0;
    int_out25 = 0;
    int_in26 = 0;
    int_out26 = 0;
    int_in27 = 0;
    int_out27 = 0;
    int_in28 = 0;
    int_out28 = 0;
    int_in29 = 0;
    int_out29 = 0;
    int_in30 = 0;
    int_out30 = 0;
    int_in31 = 0;
    int_out31 = 0;
  end


endmodule



module app_top #
(
  parameter C_M_AXI_ADDR_WIDTH = 64,
  parameter C_M_AXI_DATA_WIDTH = 256
)
(
  input ap_clk,
  input ap_rst_n,
  output m00_axi_awvalid,
  input m00_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m00_axi_awaddr,
  output [8-1:0] m00_axi_awlen,
  output m00_axi_wvalid,
  input m00_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m00_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m00_axi_wstrb,
  output m00_axi_wlast,
  input m00_axi_bvalid,
  output m00_axi_bready,
  output m00_axi_arvalid,
  input m00_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m00_axi_araddr,
  output [8-1:0] m00_axi_arlen,
  input m00_axi_rvalid,
  output m00_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m00_axi_rdata,
  input m00_axi_rlast,
  output m01_axi_awvalid,
  input m01_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m01_axi_awaddr,
  output [8-1:0] m01_axi_awlen,
  output m01_axi_wvalid,
  input m01_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m01_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m01_axi_wstrb,
  output m01_axi_wlast,
  input m01_axi_bvalid,
  output m01_axi_bready,
  output m01_axi_arvalid,
  input m01_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m01_axi_araddr,
  output [8-1:0] m01_axi_arlen,
  input m01_axi_rvalid,
  output m01_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m01_axi_rdata,
  input m01_axi_rlast,
  output m02_axi_awvalid,
  input m02_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m02_axi_awaddr,
  output [8-1:0] m02_axi_awlen,
  output m02_axi_wvalid,
  input m02_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m02_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m02_axi_wstrb,
  output m02_axi_wlast,
  input m02_axi_bvalid,
  output m02_axi_bready,
  output m02_axi_arvalid,
  input m02_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m02_axi_araddr,
  output [8-1:0] m02_axi_arlen,
  input m02_axi_rvalid,
  output m02_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m02_axi_rdata,
  input m02_axi_rlast,
  output m03_axi_awvalid,
  input m03_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m03_axi_awaddr,
  output [8-1:0] m03_axi_awlen,
  output m03_axi_wvalid,
  input m03_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m03_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m03_axi_wstrb,
  output m03_axi_wlast,
  input m03_axi_bvalid,
  output m03_axi_bready,
  output m03_axi_arvalid,
  input m03_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m03_axi_araddr,
  output [8-1:0] m03_axi_arlen,
  input m03_axi_rvalid,
  output m03_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m03_axi_rdata,
  input m03_axi_rlast,
  output m04_axi_awvalid,
  input m04_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m04_axi_awaddr,
  output [8-1:0] m04_axi_awlen,
  output m04_axi_wvalid,
  input m04_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m04_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m04_axi_wstrb,
  output m04_axi_wlast,
  input m04_axi_bvalid,
  output m04_axi_bready,
  output m04_axi_arvalid,
  input m04_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m04_axi_araddr,
  output [8-1:0] m04_axi_arlen,
  input m04_axi_rvalid,
  output m04_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m04_axi_rdata,
  input m04_axi_rlast,
  output m05_axi_awvalid,
  input m05_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m05_axi_awaddr,
  output [8-1:0] m05_axi_awlen,
  output m05_axi_wvalid,
  input m05_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m05_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m05_axi_wstrb,
  output m05_axi_wlast,
  input m05_axi_bvalid,
  output m05_axi_bready,
  output m05_axi_arvalid,
  input m05_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m05_axi_araddr,
  output [8-1:0] m05_axi_arlen,
  input m05_axi_rvalid,
  output m05_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m05_axi_rdata,
  input m05_axi_rlast,
  output m06_axi_awvalid,
  input m06_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m06_axi_awaddr,
  output [8-1:0] m06_axi_awlen,
  output m06_axi_wvalid,
  input m06_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m06_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m06_axi_wstrb,
  output m06_axi_wlast,
  input m06_axi_bvalid,
  output m06_axi_bready,
  output m06_axi_arvalid,
  input m06_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m06_axi_araddr,
  output [8-1:0] m06_axi_arlen,
  input m06_axi_rvalid,
  output m06_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m06_axi_rdata,
  input m06_axi_rlast,
  output m07_axi_awvalid,
  input m07_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m07_axi_awaddr,
  output [8-1:0] m07_axi_awlen,
  output m07_axi_wvalid,
  input m07_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m07_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m07_axi_wstrb,
  output m07_axi_wlast,
  input m07_axi_bvalid,
  output m07_axi_bready,
  output m07_axi_arvalid,
  input m07_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m07_axi_araddr,
  output [8-1:0] m07_axi_arlen,
  input m07_axi_rvalid,
  output m07_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m07_axi_rdata,
  input m07_axi_rlast,
  output m08_axi_awvalid,
  input m08_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m08_axi_awaddr,
  output [8-1:0] m08_axi_awlen,
  output m08_axi_wvalid,
  input m08_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m08_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m08_axi_wstrb,
  output m08_axi_wlast,
  input m08_axi_bvalid,
  output m08_axi_bready,
  output m08_axi_arvalid,
  input m08_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m08_axi_araddr,
  output [8-1:0] m08_axi_arlen,
  input m08_axi_rvalid,
  output m08_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m08_axi_rdata,
  input m08_axi_rlast,
  output m09_axi_awvalid,
  input m09_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m09_axi_awaddr,
  output [8-1:0] m09_axi_awlen,
  output m09_axi_wvalid,
  input m09_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m09_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m09_axi_wstrb,
  output m09_axi_wlast,
  input m09_axi_bvalid,
  output m09_axi_bready,
  output m09_axi_arvalid,
  input m09_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m09_axi_araddr,
  output [8-1:0] m09_axi_arlen,
  input m09_axi_rvalid,
  output m09_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m09_axi_rdata,
  input m09_axi_rlast,
  output m10_axi_awvalid,
  input m10_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m10_axi_awaddr,
  output [8-1:0] m10_axi_awlen,
  output m10_axi_wvalid,
  input m10_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m10_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m10_axi_wstrb,
  output m10_axi_wlast,
  input m10_axi_bvalid,
  output m10_axi_bready,
  output m10_axi_arvalid,
  input m10_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m10_axi_araddr,
  output [8-1:0] m10_axi_arlen,
  input m10_axi_rvalid,
  output m10_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m10_axi_rdata,
  input m10_axi_rlast,
  output m11_axi_awvalid,
  input m11_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m11_axi_awaddr,
  output [8-1:0] m11_axi_awlen,
  output m11_axi_wvalid,
  input m11_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m11_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m11_axi_wstrb,
  output m11_axi_wlast,
  input m11_axi_bvalid,
  output m11_axi_bready,
  output m11_axi_arvalid,
  input m11_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m11_axi_araddr,
  output [8-1:0] m11_axi_arlen,
  input m11_axi_rvalid,
  output m11_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m11_axi_rdata,
  input m11_axi_rlast,
  output m12_axi_awvalid,
  input m12_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m12_axi_awaddr,
  output [8-1:0] m12_axi_awlen,
  output m12_axi_wvalid,
  input m12_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m12_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m12_axi_wstrb,
  output m12_axi_wlast,
  input m12_axi_bvalid,
  output m12_axi_bready,
  output m12_axi_arvalid,
  input m12_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m12_axi_araddr,
  output [8-1:0] m12_axi_arlen,
  input m12_axi_rvalid,
  output m12_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m12_axi_rdata,
  input m12_axi_rlast,
  output m13_axi_awvalid,
  input m13_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m13_axi_awaddr,
  output [8-1:0] m13_axi_awlen,
  output m13_axi_wvalid,
  input m13_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m13_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m13_axi_wstrb,
  output m13_axi_wlast,
  input m13_axi_bvalid,
  output m13_axi_bready,
  output m13_axi_arvalid,
  input m13_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m13_axi_araddr,
  output [8-1:0] m13_axi_arlen,
  input m13_axi_rvalid,
  output m13_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m13_axi_rdata,
  input m13_axi_rlast,
  output m14_axi_awvalid,
  input m14_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m14_axi_awaddr,
  output [8-1:0] m14_axi_awlen,
  output m14_axi_wvalid,
  input m14_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m14_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m14_axi_wstrb,
  output m14_axi_wlast,
  input m14_axi_bvalid,
  output m14_axi_bready,
  output m14_axi_arvalid,
  input m14_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m14_axi_araddr,
  output [8-1:0] m14_axi_arlen,
  input m14_axi_rvalid,
  output m14_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m14_axi_rdata,
  input m14_axi_rlast,
  output m15_axi_awvalid,
  input m15_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m15_axi_awaddr,
  output [8-1:0] m15_axi_awlen,
  output m15_axi_wvalid,
  input m15_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m15_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m15_axi_wstrb,
  output m15_axi_wlast,
  input m15_axi_bvalid,
  output m15_axi_bready,
  output m15_axi_arvalid,
  input m15_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m15_axi_araddr,
  output [8-1:0] m15_axi_arlen,
  input m15_axi_rvalid,
  output m15_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m15_axi_rdata,
  input m15_axi_rlast,
  output m16_axi_awvalid,
  input m16_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m16_axi_awaddr,
  output [8-1:0] m16_axi_awlen,
  output m16_axi_wvalid,
  input m16_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m16_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m16_axi_wstrb,
  output m16_axi_wlast,
  input m16_axi_bvalid,
  output m16_axi_bready,
  output m16_axi_arvalid,
  input m16_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m16_axi_araddr,
  output [8-1:0] m16_axi_arlen,
  input m16_axi_rvalid,
  output m16_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m16_axi_rdata,
  input m16_axi_rlast,
  output m17_axi_awvalid,
  input m17_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m17_axi_awaddr,
  output [8-1:0] m17_axi_awlen,
  output m17_axi_wvalid,
  input m17_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m17_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m17_axi_wstrb,
  output m17_axi_wlast,
  input m17_axi_bvalid,
  output m17_axi_bready,
  output m17_axi_arvalid,
  input m17_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m17_axi_araddr,
  output [8-1:0] m17_axi_arlen,
  input m17_axi_rvalid,
  output m17_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m17_axi_rdata,
  input m17_axi_rlast,
  output m18_axi_awvalid,
  input m18_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m18_axi_awaddr,
  output [8-1:0] m18_axi_awlen,
  output m18_axi_wvalid,
  input m18_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m18_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m18_axi_wstrb,
  output m18_axi_wlast,
  input m18_axi_bvalid,
  output m18_axi_bready,
  output m18_axi_arvalid,
  input m18_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m18_axi_araddr,
  output [8-1:0] m18_axi_arlen,
  input m18_axi_rvalid,
  output m18_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m18_axi_rdata,
  input m18_axi_rlast,
  output m19_axi_awvalid,
  input m19_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m19_axi_awaddr,
  output [8-1:0] m19_axi_awlen,
  output m19_axi_wvalid,
  input m19_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m19_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m19_axi_wstrb,
  output m19_axi_wlast,
  input m19_axi_bvalid,
  output m19_axi_bready,
  output m19_axi_arvalid,
  input m19_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m19_axi_araddr,
  output [8-1:0] m19_axi_arlen,
  input m19_axi_rvalid,
  output m19_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m19_axi_rdata,
  input m19_axi_rlast,
  output m20_axi_awvalid,
  input m20_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m20_axi_awaddr,
  output [8-1:0] m20_axi_awlen,
  output m20_axi_wvalid,
  input m20_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m20_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m20_axi_wstrb,
  output m20_axi_wlast,
  input m20_axi_bvalid,
  output m20_axi_bready,
  output m20_axi_arvalid,
  input m20_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m20_axi_araddr,
  output [8-1:0] m20_axi_arlen,
  input m20_axi_rvalid,
  output m20_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m20_axi_rdata,
  input m20_axi_rlast,
  output m21_axi_awvalid,
  input m21_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m21_axi_awaddr,
  output [8-1:0] m21_axi_awlen,
  output m21_axi_wvalid,
  input m21_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m21_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m21_axi_wstrb,
  output m21_axi_wlast,
  input m21_axi_bvalid,
  output m21_axi_bready,
  output m21_axi_arvalid,
  input m21_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m21_axi_araddr,
  output [8-1:0] m21_axi_arlen,
  input m21_axi_rvalid,
  output m21_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m21_axi_rdata,
  input m21_axi_rlast,
  output m22_axi_awvalid,
  input m22_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m22_axi_awaddr,
  output [8-1:0] m22_axi_awlen,
  output m22_axi_wvalid,
  input m22_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m22_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m22_axi_wstrb,
  output m22_axi_wlast,
  input m22_axi_bvalid,
  output m22_axi_bready,
  output m22_axi_arvalid,
  input m22_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m22_axi_araddr,
  output [8-1:0] m22_axi_arlen,
  input m22_axi_rvalid,
  output m22_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m22_axi_rdata,
  input m22_axi_rlast,
  output m23_axi_awvalid,
  input m23_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m23_axi_awaddr,
  output [8-1:0] m23_axi_awlen,
  output m23_axi_wvalid,
  input m23_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m23_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m23_axi_wstrb,
  output m23_axi_wlast,
  input m23_axi_bvalid,
  output m23_axi_bready,
  output m23_axi_arvalid,
  input m23_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m23_axi_araddr,
  output [8-1:0] m23_axi_arlen,
  input m23_axi_rvalid,
  output m23_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m23_axi_rdata,
  input m23_axi_rlast,
  output m24_axi_awvalid,
  input m24_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m24_axi_awaddr,
  output [8-1:0] m24_axi_awlen,
  output m24_axi_wvalid,
  input m24_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m24_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m24_axi_wstrb,
  output m24_axi_wlast,
  input m24_axi_bvalid,
  output m24_axi_bready,
  output m24_axi_arvalid,
  input m24_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m24_axi_araddr,
  output [8-1:0] m24_axi_arlen,
  input m24_axi_rvalid,
  output m24_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m24_axi_rdata,
  input m24_axi_rlast,
  output m25_axi_awvalid,
  input m25_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m25_axi_awaddr,
  output [8-1:0] m25_axi_awlen,
  output m25_axi_wvalid,
  input m25_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m25_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m25_axi_wstrb,
  output m25_axi_wlast,
  input m25_axi_bvalid,
  output m25_axi_bready,
  output m25_axi_arvalid,
  input m25_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m25_axi_araddr,
  output [8-1:0] m25_axi_arlen,
  input m25_axi_rvalid,
  output m25_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m25_axi_rdata,
  input m25_axi_rlast,
  output m26_axi_awvalid,
  input m26_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m26_axi_awaddr,
  output [8-1:0] m26_axi_awlen,
  output m26_axi_wvalid,
  input m26_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m26_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m26_axi_wstrb,
  output m26_axi_wlast,
  input m26_axi_bvalid,
  output m26_axi_bready,
  output m26_axi_arvalid,
  input m26_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m26_axi_araddr,
  output [8-1:0] m26_axi_arlen,
  input m26_axi_rvalid,
  output m26_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m26_axi_rdata,
  input m26_axi_rlast,
  output m27_axi_awvalid,
  input m27_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m27_axi_awaddr,
  output [8-1:0] m27_axi_awlen,
  output m27_axi_wvalid,
  input m27_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m27_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m27_axi_wstrb,
  output m27_axi_wlast,
  input m27_axi_bvalid,
  output m27_axi_bready,
  output m27_axi_arvalid,
  input m27_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m27_axi_araddr,
  output [8-1:0] m27_axi_arlen,
  input m27_axi_rvalid,
  output m27_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m27_axi_rdata,
  input m27_axi_rlast,
  output m28_axi_awvalid,
  input m28_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m28_axi_awaddr,
  output [8-1:0] m28_axi_awlen,
  output m28_axi_wvalid,
  input m28_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m28_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m28_axi_wstrb,
  output m28_axi_wlast,
  input m28_axi_bvalid,
  output m28_axi_bready,
  output m28_axi_arvalid,
  input m28_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m28_axi_araddr,
  output [8-1:0] m28_axi_arlen,
  input m28_axi_rvalid,
  output m28_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m28_axi_rdata,
  input m28_axi_rlast,
  output m29_axi_awvalid,
  input m29_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m29_axi_awaddr,
  output [8-1:0] m29_axi_awlen,
  output m29_axi_wvalid,
  input m29_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m29_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m29_axi_wstrb,
  output m29_axi_wlast,
  input m29_axi_bvalid,
  output m29_axi_bready,
  output m29_axi_arvalid,
  input m29_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m29_axi_araddr,
  output [8-1:0] m29_axi_arlen,
  input m29_axi_rvalid,
  output m29_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m29_axi_rdata,
  input m29_axi_rlast,
  output m30_axi_awvalid,
  input m30_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m30_axi_awaddr,
  output [8-1:0] m30_axi_awlen,
  output m30_axi_wvalid,
  input m30_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m30_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m30_axi_wstrb,
  output m30_axi_wlast,
  input m30_axi_bvalid,
  output m30_axi_bready,
  output m30_axi_arvalid,
  input m30_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m30_axi_araddr,
  output [8-1:0] m30_axi_arlen,
  input m30_axi_rvalid,
  output m30_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m30_axi_rdata,
  input m30_axi_rlast,
  output m31_axi_awvalid,
  input m31_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m31_axi_awaddr,
  output [8-1:0] m31_axi_awlen,
  output m31_axi_wvalid,
  input m31_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m31_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m31_axi_wstrb,
  output m31_axi_wlast,
  input m31_axi_bvalid,
  output m31_axi_bready,
  output m31_axi_arvalid,
  input m31_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m31_axi_araddr,
  output [8-1:0] m31_axi_arlen,
  input m31_axi_rvalid,
  output m31_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m31_axi_rdata,
  input m31_axi_rlast,
  input ap_start,
  output ap_idle,
  output ap_done,
  output ap_ready,
  input [32-1:0] in_s0,
  input [32-1:0] in_s1,
  input [32-1:0] in_s2,
  input [32-1:0] in_s3,
  input [32-1:0] in_s4,
  input [32-1:0] in_s5,
  input [32-1:0] in_s6,
  input [32-1:0] in_s7,
  input [32-1:0] in_s8,
  input [32-1:0] in_s9,
  input [32-1:0] in_s10,
  input [32-1:0] in_s11,
  input [32-1:0] in_s12,
  input [32-1:0] in_s13,
  input [32-1:0] in_s14,
  input [32-1:0] in_s15,
  input [32-1:0] in_s16,
  input [32-1:0] in_s17,
  input [32-1:0] in_s18,
  input [32-1:0] in_s19,
  input [32-1:0] in_s20,
  input [32-1:0] in_s21,
  input [32-1:0] in_s22,
  input [32-1:0] in_s23,
  input [32-1:0] in_s24,
  input [32-1:0] in_s25,
  input [32-1:0] in_s26,
  input [32-1:0] in_s27,
  input [32-1:0] in_s28,
  input [32-1:0] in_s29,
  input [32-1:0] in_s30,
  input [32-1:0] in_s31,
  input [32-1:0] out_s0,
  input [32-1:0] out_s1,
  input [32-1:0] out_s2,
  input [32-1:0] out_s3,
  input [32-1:0] out_s4,
  input [32-1:0] out_s5,
  input [32-1:0] out_s6,
  input [32-1:0] out_s7,
  input [32-1:0] out_s8,
  input [32-1:0] out_s9,
  input [32-1:0] out_s10,
  input [32-1:0] out_s11,
  input [32-1:0] out_s12,
  input [32-1:0] out_s13,
  input [32-1:0] out_s14,
  input [32-1:0] out_s15,
  input [32-1:0] out_s16,
  input [32-1:0] out_s17,
  input [32-1:0] out_s18,
  input [32-1:0] out_s19,
  input [32-1:0] out_s20,
  input [32-1:0] out_s21,
  input [32-1:0] out_s22,
  input [32-1:0] out_s23,
  input [32-1:0] out_s24,
  input [32-1:0] out_s25,
  input [32-1:0] out_s26,
  input [32-1:0] out_s27,
  input [32-1:0] out_s28,
  input [32-1:0] out_s29,
  input [32-1:0] out_s30,
  input [32-1:0] out_s31,
  input [64-1:0] in0,
  input [64-1:0] out0,
  input [64-1:0] in1,
  input [64-1:0] out1,
  input [64-1:0] in2,
  input [64-1:0] out2,
  input [64-1:0] in3,
  input [64-1:0] out3,
  input [64-1:0] in4,
  input [64-1:0] out4,
  input [64-1:0] in5,
  input [64-1:0] out5,
  input [64-1:0] in6,
  input [64-1:0] out6,
  input [64-1:0] in7,
  input [64-1:0] out7,
  input [64-1:0] in8,
  input [64-1:0] out8,
  input [64-1:0] in9,
  input [64-1:0] out9,
  input [64-1:0] in10,
  input [64-1:0] out10,
  input [64-1:0] in11,
  input [64-1:0] out11,
  input [64-1:0] in12,
  input [64-1:0] out12,
  input [64-1:0] in13,
  input [64-1:0] out13,
  input [64-1:0] in14,
  input [64-1:0] out14,
  input [64-1:0] in15,
  input [64-1:0] out15,
  input [64-1:0] in16,
  input [64-1:0] out16,
  input [64-1:0] in17,
  input [64-1:0] out17,
  input [64-1:0] in18,
  input [64-1:0] out18,
  input [64-1:0] in19,
  input [64-1:0] out19,
  input [64-1:0] in20,
  input [64-1:0] out20,
  input [64-1:0] in21,
  input [64-1:0] out21,
  input [64-1:0] in22,
  input [64-1:0] out22,
  input [64-1:0] in23,
  input [64-1:0] out23,
  input [64-1:0] in24,
  input [64-1:0] out24,
  input [64-1:0] in25,
  input [64-1:0] out25,
  input [64-1:0] in26,
  input [64-1:0] out26,
  input [64-1:0] in27,
  input [64-1:0] out27,
  input [64-1:0] in28,
  input [64-1:0] out28,
  input [64-1:0] in29,
  input [64-1:0] out29,
  input [64-1:0] in30,
  input [64-1:0] out30,
  input [64-1:0] in31,
  input [64-1:0] out31
);

  localparam LP_NUM_EXAMPLES = 32;
  localparam LP_RD_MAX_OUTSTANDING = 16;
  localparam LP_WR_MAX_OUTSTANDING = 16;
  (* KEEP = "yes" *)
  reg reset;
  reg ap_idle_r;
  reg ap_done_r;
  wire [LP_NUM_EXAMPLES-1:0] rd_ctrl_done;
  wire [LP_NUM_EXAMPLES-1:0] wr_ctrl_done;
  reg [LP_NUM_EXAMPLES-1:0] acc_user_done_rd_data;
  reg [LP_NUM_EXAMPLES-1:0] acc_user_done_wr_data;
  wire [LP_NUM_EXAMPLES-1:0] acc_user_request_read;
  wire [LP_NUM_EXAMPLES-1:0] acc_user_read_data_valid;
  wire [C_M_AXI_DATA_WIDTH*LP_NUM_EXAMPLES-1:0] acc_user_read_data;
  wire [LP_NUM_EXAMPLES-1:0] acc_user_available_write;
  wire [LP_NUM_EXAMPLES-1:0] acc_user_request_write;
  wire [C_M_AXI_DATA_WIDTH*LP_NUM_EXAMPLES-1:0] acc_user_write_data;
  wire acc_user_done;
  wire rd_tvalid0;
  wire rd_tready0;
  wire rd_tlast0;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata0;
  wire rd_tvalid1;
  wire rd_tready1;
  wire rd_tlast1;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata1;
  wire rd_tvalid2;
  wire rd_tready2;
  wire rd_tlast2;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata2;
  wire rd_tvalid3;
  wire rd_tready3;
  wire rd_tlast3;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata3;
  wire rd_tvalid4;
  wire rd_tready4;
  wire rd_tlast4;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata4;
  wire rd_tvalid5;
  wire rd_tready5;
  wire rd_tlast5;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata5;
  wire rd_tvalid6;
  wire rd_tready6;
  wire rd_tlast6;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata6;
  wire rd_tvalid7;
  wire rd_tready7;
  wire rd_tlast7;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata7;
  wire rd_tvalid8;
  wire rd_tready8;
  wire rd_tlast8;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata8;
  wire rd_tvalid9;
  wire rd_tready9;
  wire rd_tlast9;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata9;
  wire rd_tvalid10;
  wire rd_tready10;
  wire rd_tlast10;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata10;
  wire rd_tvalid11;
  wire rd_tready11;
  wire rd_tlast11;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata11;
  wire rd_tvalid12;
  wire rd_tready12;
  wire rd_tlast12;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata12;
  wire rd_tvalid13;
  wire rd_tready13;
  wire rd_tlast13;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata13;
  wire rd_tvalid14;
  wire rd_tready14;
  wire rd_tlast14;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata14;
  wire rd_tvalid15;
  wire rd_tready15;
  wire rd_tlast15;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata15;
  wire rd_tvalid16;
  wire rd_tready16;
  wire rd_tlast16;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata16;
  wire rd_tvalid17;
  wire rd_tready17;
  wire rd_tlast17;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata17;
  wire rd_tvalid18;
  wire rd_tready18;
  wire rd_tlast18;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata18;
  wire rd_tvalid19;
  wire rd_tready19;
  wire rd_tlast19;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata19;
  wire rd_tvalid20;
  wire rd_tready20;
  wire rd_tlast20;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata20;
  wire rd_tvalid21;
  wire rd_tready21;
  wire rd_tlast21;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata21;
  wire rd_tvalid22;
  wire rd_tready22;
  wire rd_tlast22;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata22;
  wire rd_tvalid23;
  wire rd_tready23;
  wire rd_tlast23;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata23;
  wire rd_tvalid24;
  wire rd_tready24;
  wire rd_tlast24;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata24;
  wire rd_tvalid25;
  wire rd_tready25;
  wire rd_tlast25;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata25;
  wire rd_tvalid26;
  wire rd_tready26;
  wire rd_tlast26;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata26;
  wire rd_tvalid27;
  wire rd_tready27;
  wire rd_tlast27;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata27;
  wire rd_tvalid28;
  wire rd_tready28;
  wire rd_tlast28;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata28;
  wire rd_tvalid29;
  wire rd_tready29;
  wire rd_tlast29;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata29;
  wire rd_tvalid30;
  wire rd_tready30;
  wire rd_tlast30;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata30;
  wire rd_tvalid31;
  wire rd_tready31;
  wire rd_tlast31;
  wire [C_M_AXI_DATA_WIDTH-1:0] rd_tdata31;
  wire wr_tvalid0;
  wire wr_tready0;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata0;
  wire wr_tvalid1;
  wire wr_tready1;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata1;
  wire wr_tvalid2;
  wire wr_tready2;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata2;
  wire wr_tvalid3;
  wire wr_tready3;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata3;
  wire wr_tvalid4;
  wire wr_tready4;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata4;
  wire wr_tvalid5;
  wire wr_tready5;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata5;
  wire wr_tvalid6;
  wire wr_tready6;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata6;
  wire wr_tvalid7;
  wire wr_tready7;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata7;
  wire wr_tvalid8;
  wire wr_tready8;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata8;
  wire wr_tvalid9;
  wire wr_tready9;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata9;
  wire wr_tvalid10;
  wire wr_tready10;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata10;
  wire wr_tvalid11;
  wire wr_tready11;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata11;
  wire wr_tvalid12;
  wire wr_tready12;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata12;
  wire wr_tvalid13;
  wire wr_tready13;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata13;
  wire wr_tvalid14;
  wire wr_tready14;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata14;
  wire wr_tvalid15;
  wire wr_tready15;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata15;
  wire wr_tvalid16;
  wire wr_tready16;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata16;
  wire wr_tvalid17;
  wire wr_tready17;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata17;
  wire wr_tvalid18;
  wire wr_tready18;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata18;
  wire wr_tvalid19;
  wire wr_tready19;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata19;
  wire wr_tvalid20;
  wire wr_tready20;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata20;
  wire wr_tvalid21;
  wire wr_tready21;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata21;
  wire wr_tvalid22;
  wire wr_tready22;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata22;
  wire wr_tvalid23;
  wire wr_tready23;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata23;
  wire wr_tvalid24;
  wire wr_tready24;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata24;
  wire wr_tvalid25;
  wire wr_tready25;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata25;
  wire wr_tvalid26;
  wire wr_tready26;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata26;
  wire wr_tvalid27;
  wire wr_tready27;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata27;
  wire wr_tvalid28;
  wire wr_tready28;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata28;
  wire wr_tvalid29;
  wire wr_tready29;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata29;
  wire wr_tvalid30;
  wire wr_tready30;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata30;
  wire wr_tvalid31;
  wire wr_tready31;
  wire [C_M_AXI_DATA_WIDTH-1:0] wr_tdata31;
  reg [2-1:0] fsm_reset;
  reg areset;
  reg ap_start_pulse;
  reg user_start;
  localparam FSM_STATE_START = 2'b0;
  localparam FSM_STATE_RESET = 2'b1;
  localparam FSM_STATE_RUNNING = 2'b10;

  always @(posedge ap_clk) begin
    reset <= ~ap_rst_n;
  end


  always @(posedge ap_clk) begin
    if(reset) begin
      areset <= 1'b0;
      fsm_reset <= FSM_STATE_START;
      ap_start_pulse <= 1'b0;
      user_start <= 1'b0;
    end else begin
      areset <= 1'b0;
      ap_start_pulse <= 1'b0;
      case(fsm_reset)
        FSM_STATE_START: begin
          if(ap_start) begin
            areset <= 1'b1;
            fsm_reset <= FSM_STATE_RESET;
            user_start <= 1'b0;
          end 
        end
        FSM_STATE_RESET: begin
          ap_start_pulse <= 1'b1;
          user_start <= 1'b1;
          fsm_reset <= FSM_STATE_RUNNING;
        end
        FSM_STATE_RUNNING: begin
          if(~ap_start) begin
            fsm_reset <= FSM_STATE_START;
          end 
        end
      endcase
    end
  end


  always @(posedge ap_clk) begin
    if(areset) begin
      ap_idle_r <= 1'b1;
    end else begin
      ap_idle_r <= (ap_done)? 1'b1 : 
                   (ap_start_pulse)? 1'b0 : ap_idle;
    end
  end

  assign ap_idle = ap_idle_r;

  always @(posedge ap_clk) begin
    if(areset) begin
      ap_done_r <= 1'b0;
    end else begin
      ap_done_r <= (ap_done)? 1'b0 : ap_done_r | acc_user_done;
    end
  end

  assign ap_done = ap_done_r;
  assign ap_ready = ap_done;
  integer i;

  always @(posedge ap_clk) begin
    if(areset) begin
      acc_user_done_rd_data <= { LP_NUM_EXAMPLES{ 1'b0 } };
      acc_user_done_wr_data <= { LP_NUM_EXAMPLES{ 1'b0 } };
    end else begin
      for(i=0; i<LP_NUM_EXAMPLES; i=i+1) begin
        acc_user_done_rd_data[i] <= (rd_ctrl_done[i])? 1'b1 : acc_user_done_rd_data[i];
        acc_user_done_wr_data[i] <= (wr_ctrl_done[i])? 1'b1 : acc_user_done_wr_data[i];
      end
    end
  end

  assign rd_tready0 = acc_user_request_read[0];
  assign rd_tready1 = acc_user_request_read[1];
  assign rd_tready2 = acc_user_request_read[2];
  assign rd_tready3 = acc_user_request_read[3];
  assign rd_tready4 = acc_user_request_read[4];
  assign rd_tready5 = acc_user_request_read[5];
  assign rd_tready6 = acc_user_request_read[6];
  assign rd_tready7 = acc_user_request_read[7];
  assign rd_tready8 = acc_user_request_read[8];
  assign rd_tready9 = acc_user_request_read[9];
  assign rd_tready10 = acc_user_request_read[10];
  assign rd_tready11 = acc_user_request_read[11];
  assign rd_tready12 = acc_user_request_read[12];
  assign rd_tready13 = acc_user_request_read[13];
  assign rd_tready14 = acc_user_request_read[14];
  assign rd_tready15 = acc_user_request_read[15];
  assign rd_tready16 = acc_user_request_read[16];
  assign rd_tready17 = acc_user_request_read[17];
  assign rd_tready18 = acc_user_request_read[18];
  assign rd_tready19 = acc_user_request_read[19];
  assign rd_tready20 = acc_user_request_read[20];
  assign rd_tready21 = acc_user_request_read[21];
  assign rd_tready22 = acc_user_request_read[22];
  assign rd_tready23 = acc_user_request_read[23];
  assign rd_tready24 = acc_user_request_read[24];
  assign rd_tready25 = acc_user_request_read[25];
  assign rd_tready26 = acc_user_request_read[26];
  assign rd_tready27 = acc_user_request_read[27];
  assign rd_tready28 = acc_user_request_read[28];
  assign rd_tready29 = acc_user_request_read[29];
  assign rd_tready30 = acc_user_request_read[30];
  assign rd_tready31 = acc_user_request_read[31];
  assign acc_user_read_data_valid = {rd_tvalid31,rd_tvalid30,rd_tvalid29,rd_tvalid28,rd_tvalid27,rd_tvalid26,rd_tvalid25,rd_tvalid24,rd_tvalid23,rd_tvalid22,rd_tvalid21,rd_tvalid20,rd_tvalid19,rd_tvalid18,rd_tvalid17,rd_tvalid16,rd_tvalid15,rd_tvalid14,rd_tvalid13,rd_tvalid12,rd_tvalid11,rd_tvalid10,rd_tvalid9,rd_tvalid8,rd_tvalid7,rd_tvalid6,rd_tvalid5,rd_tvalid4,rd_tvalid3,rd_tvalid2,rd_tvalid1,rd_tvalid0};
  assign acc_user_read_data = {rd_tdata31,rd_tdata30,rd_tdata29,rd_tdata28,rd_tdata27,rd_tdata26,rd_tdata25,rd_tdata24,rd_tdata23,rd_tdata22,rd_tdata21,rd_tdata20,rd_tdata19,rd_tdata18,rd_tdata17,rd_tdata16,rd_tdata15,rd_tdata14,rd_tdata13,rd_tdata12,rd_tdata11,rd_tdata10,rd_tdata9,rd_tdata8,rd_tdata7,rd_tdata6,rd_tdata5,rd_tdata4,rd_tdata3,rd_tdata2,rd_tdata1,rd_tdata0};

  assign acc_user_available_write = {wr_tready31,wr_tready30,wr_tready29,wr_tready28,wr_tready27,wr_tready26,wr_tready25,wr_tready24,wr_tready23,wr_tready22,wr_tready21,wr_tready20,wr_tready19,wr_tready18,wr_tready17,wr_tready16,wr_tready15,wr_tready14,wr_tready13,wr_tready12,wr_tready11,wr_tready10,wr_tready9,wr_tready8,wr_tready7,wr_tready6,wr_tready5,wr_tready4,wr_tready3,wr_tready2,wr_tready1,wr_tready0};
  assign wr_tvalid0 = acc_user_request_write[0];
  assign wr_tdata0 = acc_user_write_data[1*C_M_AXI_DATA_WIDTH-1:0*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid1 = acc_user_request_write[1];
  assign wr_tdata1 = acc_user_write_data[2*C_M_AXI_DATA_WIDTH-1:1*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid2 = acc_user_request_write[2];
  assign wr_tdata2 = acc_user_write_data[3*C_M_AXI_DATA_WIDTH-1:2*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid3 = acc_user_request_write[3];
  assign wr_tdata3 = acc_user_write_data[4*C_M_AXI_DATA_WIDTH-1:3*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid4 = acc_user_request_write[4];
  assign wr_tdata4 = acc_user_write_data[5*C_M_AXI_DATA_WIDTH-1:4*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid5 = acc_user_request_write[5];
  assign wr_tdata5 = acc_user_write_data[6*C_M_AXI_DATA_WIDTH-1:5*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid6 = acc_user_request_write[6];
  assign wr_tdata6 = acc_user_write_data[7*C_M_AXI_DATA_WIDTH-1:6*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid7 = acc_user_request_write[7];
  assign wr_tdata7 = acc_user_write_data[8*C_M_AXI_DATA_WIDTH-1:7*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid8 = acc_user_request_write[8];
  assign wr_tdata8 = acc_user_write_data[9*C_M_AXI_DATA_WIDTH-1:8*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid9 = acc_user_request_write[9];
  assign wr_tdata9 = acc_user_write_data[10*C_M_AXI_DATA_WIDTH-1:9*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid10 = acc_user_request_write[10];
  assign wr_tdata10 = acc_user_write_data[11*C_M_AXI_DATA_WIDTH-1:10*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid11 = acc_user_request_write[11];
  assign wr_tdata11 = acc_user_write_data[12*C_M_AXI_DATA_WIDTH-1:11*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid12 = acc_user_request_write[12];
  assign wr_tdata12 = acc_user_write_data[13*C_M_AXI_DATA_WIDTH-1:12*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid13 = acc_user_request_write[13];
  assign wr_tdata13 = acc_user_write_data[14*C_M_AXI_DATA_WIDTH-1:13*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid14 = acc_user_request_write[14];
  assign wr_tdata14 = acc_user_write_data[15*C_M_AXI_DATA_WIDTH-1:14*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid15 = acc_user_request_write[15];
  assign wr_tdata15 = acc_user_write_data[16*C_M_AXI_DATA_WIDTH-1:15*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid16 = acc_user_request_write[16];
  assign wr_tdata16 = acc_user_write_data[17*C_M_AXI_DATA_WIDTH-1:16*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid17 = acc_user_request_write[17];
  assign wr_tdata17 = acc_user_write_data[18*C_M_AXI_DATA_WIDTH-1:17*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid18 = acc_user_request_write[18];
  assign wr_tdata18 = acc_user_write_data[19*C_M_AXI_DATA_WIDTH-1:18*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid19 = acc_user_request_write[19];
  assign wr_tdata19 = acc_user_write_data[20*C_M_AXI_DATA_WIDTH-1:19*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid20 = acc_user_request_write[20];
  assign wr_tdata20 = acc_user_write_data[21*C_M_AXI_DATA_WIDTH-1:20*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid21 = acc_user_request_write[21];
  assign wr_tdata21 = acc_user_write_data[22*C_M_AXI_DATA_WIDTH-1:21*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid22 = acc_user_request_write[22];
  assign wr_tdata22 = acc_user_write_data[23*C_M_AXI_DATA_WIDTH-1:22*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid23 = acc_user_request_write[23];
  assign wr_tdata23 = acc_user_write_data[24*C_M_AXI_DATA_WIDTH-1:23*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid24 = acc_user_request_write[24];
  assign wr_tdata24 = acc_user_write_data[25*C_M_AXI_DATA_WIDTH-1:24*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid25 = acc_user_request_write[25];
  assign wr_tdata25 = acc_user_write_data[26*C_M_AXI_DATA_WIDTH-1:25*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid26 = acc_user_request_write[26];
  assign wr_tdata26 = acc_user_write_data[27*C_M_AXI_DATA_WIDTH-1:26*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid27 = acc_user_request_write[27];
  assign wr_tdata27 = acc_user_write_data[28*C_M_AXI_DATA_WIDTH-1:27*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid28 = acc_user_request_write[28];
  assign wr_tdata28 = acc_user_write_data[29*C_M_AXI_DATA_WIDTH-1:28*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid29 = acc_user_request_write[29];
  assign wr_tdata29 = acc_user_write_data[30*C_M_AXI_DATA_WIDTH-1:29*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid30 = acc_user_request_write[30];
  assign wr_tdata30 = acc_user_write_data[31*C_M_AXI_DATA_WIDTH-1:30*C_M_AXI_DATA_WIDTH];
  assign wr_tvalid31 = acc_user_request_write[31];
  assign wr_tdata31 = acc_user_write_data[32*C_M_AXI_DATA_WIDTH-1:31*C_M_AXI_DATA_WIDTH];

  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_0
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[0]),
    .ctrl_addr_offset(in0),
    .ctrl_xfer_size_in_bytes(in_s0),
    .m_axi_arvalid(m00_axi_arvalid),
    .m_axi_arready(m00_axi_arready),
    .m_axi_araddr(m00_axi_araddr),
    .m_axi_arlen(m00_axi_arlen),
    .m_axi_rvalid(m00_axi_rvalid),
    .m_axi_rready(m00_axi_rready),
    .m_axi_rdata(m00_axi_rdata),
    .m_axi_rlast(m00_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid0),
    .m_axis_tready(rd_tready0),
    .m_axis_tlast(rd_tlast0),
    .m_axis_tdata(rd_tdata0)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_1
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[1]),
    .ctrl_addr_offset(in1),
    .ctrl_xfer_size_in_bytes(in_s1),
    .m_axi_arvalid(m01_axi_arvalid),
    .m_axi_arready(m01_axi_arready),
    .m_axi_araddr(m01_axi_araddr),
    .m_axi_arlen(m01_axi_arlen),
    .m_axi_rvalid(m01_axi_rvalid),
    .m_axi_rready(m01_axi_rready),
    .m_axi_rdata(m01_axi_rdata),
    .m_axi_rlast(m01_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid1),
    .m_axis_tready(rd_tready1),
    .m_axis_tlast(rd_tlast1),
    .m_axis_tdata(rd_tdata1)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_2
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[2]),
    .ctrl_addr_offset(in2),
    .ctrl_xfer_size_in_bytes(in_s2),
    .m_axi_arvalid(m02_axi_arvalid),
    .m_axi_arready(m02_axi_arready),
    .m_axi_araddr(m02_axi_araddr),
    .m_axi_arlen(m02_axi_arlen),
    .m_axi_rvalid(m02_axi_rvalid),
    .m_axi_rready(m02_axi_rready),
    .m_axi_rdata(m02_axi_rdata),
    .m_axi_rlast(m02_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid2),
    .m_axis_tready(rd_tready2),
    .m_axis_tlast(rd_tlast2),
    .m_axis_tdata(rd_tdata2)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_3
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[3]),
    .ctrl_addr_offset(in3),
    .ctrl_xfer_size_in_bytes(in_s3),
    .m_axi_arvalid(m03_axi_arvalid),
    .m_axi_arready(m03_axi_arready),
    .m_axi_araddr(m03_axi_araddr),
    .m_axi_arlen(m03_axi_arlen),
    .m_axi_rvalid(m03_axi_rvalid),
    .m_axi_rready(m03_axi_rready),
    .m_axi_rdata(m03_axi_rdata),
    .m_axi_rlast(m03_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid3),
    .m_axis_tready(rd_tready3),
    .m_axis_tlast(rd_tlast3),
    .m_axis_tdata(rd_tdata3)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_4
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[4]),
    .ctrl_addr_offset(in4),
    .ctrl_xfer_size_in_bytes(in_s4),
    .m_axi_arvalid(m04_axi_arvalid),
    .m_axi_arready(m04_axi_arready),
    .m_axi_araddr(m04_axi_araddr),
    .m_axi_arlen(m04_axi_arlen),
    .m_axi_rvalid(m04_axi_rvalid),
    .m_axi_rready(m04_axi_rready),
    .m_axi_rdata(m04_axi_rdata),
    .m_axi_rlast(m04_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid4),
    .m_axis_tready(rd_tready4),
    .m_axis_tlast(rd_tlast4),
    .m_axis_tdata(rd_tdata4)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_5
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[5]),
    .ctrl_addr_offset(in5),
    .ctrl_xfer_size_in_bytes(in_s5),
    .m_axi_arvalid(m05_axi_arvalid),
    .m_axi_arready(m05_axi_arready),
    .m_axi_araddr(m05_axi_araddr),
    .m_axi_arlen(m05_axi_arlen),
    .m_axi_rvalid(m05_axi_rvalid),
    .m_axi_rready(m05_axi_rready),
    .m_axi_rdata(m05_axi_rdata),
    .m_axi_rlast(m05_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid5),
    .m_axis_tready(rd_tready5),
    .m_axis_tlast(rd_tlast5),
    .m_axis_tdata(rd_tdata5)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_6
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[6]),
    .ctrl_addr_offset(in6),
    .ctrl_xfer_size_in_bytes(in_s6),
    .m_axi_arvalid(m06_axi_arvalid),
    .m_axi_arready(m06_axi_arready),
    .m_axi_araddr(m06_axi_araddr),
    .m_axi_arlen(m06_axi_arlen),
    .m_axi_rvalid(m06_axi_rvalid),
    .m_axi_rready(m06_axi_rready),
    .m_axi_rdata(m06_axi_rdata),
    .m_axi_rlast(m06_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid6),
    .m_axis_tready(rd_tready6),
    .m_axis_tlast(rd_tlast6),
    .m_axis_tdata(rd_tdata6)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_7
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[7]),
    .ctrl_addr_offset(in7),
    .ctrl_xfer_size_in_bytes(in_s7),
    .m_axi_arvalid(m07_axi_arvalid),
    .m_axi_arready(m07_axi_arready),
    .m_axi_araddr(m07_axi_araddr),
    .m_axi_arlen(m07_axi_arlen),
    .m_axi_rvalid(m07_axi_rvalid),
    .m_axi_rready(m07_axi_rready),
    .m_axi_rdata(m07_axi_rdata),
    .m_axi_rlast(m07_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid7),
    .m_axis_tready(rd_tready7),
    .m_axis_tlast(rd_tlast7),
    .m_axis_tdata(rd_tdata7)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_8
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[8]),
    .ctrl_addr_offset(in8),
    .ctrl_xfer_size_in_bytes(in_s8),
    .m_axi_arvalid(m08_axi_arvalid),
    .m_axi_arready(m08_axi_arready),
    .m_axi_araddr(m08_axi_araddr),
    .m_axi_arlen(m08_axi_arlen),
    .m_axi_rvalid(m08_axi_rvalid),
    .m_axi_rready(m08_axi_rready),
    .m_axi_rdata(m08_axi_rdata),
    .m_axi_rlast(m08_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid8),
    .m_axis_tready(rd_tready8),
    .m_axis_tlast(rd_tlast8),
    .m_axis_tdata(rd_tdata8)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_9
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[9]),
    .ctrl_addr_offset(in9),
    .ctrl_xfer_size_in_bytes(in_s9),
    .m_axi_arvalid(m09_axi_arvalid),
    .m_axi_arready(m09_axi_arready),
    .m_axi_araddr(m09_axi_araddr),
    .m_axi_arlen(m09_axi_arlen),
    .m_axi_rvalid(m09_axi_rvalid),
    .m_axi_rready(m09_axi_rready),
    .m_axi_rdata(m09_axi_rdata),
    .m_axi_rlast(m09_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid9),
    .m_axis_tready(rd_tready9),
    .m_axis_tlast(rd_tlast9),
    .m_axis_tdata(rd_tdata9)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_10
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[10]),
    .ctrl_addr_offset(in10),
    .ctrl_xfer_size_in_bytes(in_s10),
    .m_axi_arvalid(m10_axi_arvalid),
    .m_axi_arready(m10_axi_arready),
    .m_axi_araddr(m10_axi_araddr),
    .m_axi_arlen(m10_axi_arlen),
    .m_axi_rvalid(m10_axi_rvalid),
    .m_axi_rready(m10_axi_rready),
    .m_axi_rdata(m10_axi_rdata),
    .m_axi_rlast(m10_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid10),
    .m_axis_tready(rd_tready10),
    .m_axis_tlast(rd_tlast10),
    .m_axis_tdata(rd_tdata10)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_11
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[11]),
    .ctrl_addr_offset(in11),
    .ctrl_xfer_size_in_bytes(in_s11),
    .m_axi_arvalid(m11_axi_arvalid),
    .m_axi_arready(m11_axi_arready),
    .m_axi_araddr(m11_axi_araddr),
    .m_axi_arlen(m11_axi_arlen),
    .m_axi_rvalid(m11_axi_rvalid),
    .m_axi_rready(m11_axi_rready),
    .m_axi_rdata(m11_axi_rdata),
    .m_axi_rlast(m11_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid11),
    .m_axis_tready(rd_tready11),
    .m_axis_tlast(rd_tlast11),
    .m_axis_tdata(rd_tdata11)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_12
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[12]),
    .ctrl_addr_offset(in12),
    .ctrl_xfer_size_in_bytes(in_s12),
    .m_axi_arvalid(m12_axi_arvalid),
    .m_axi_arready(m12_axi_arready),
    .m_axi_araddr(m12_axi_araddr),
    .m_axi_arlen(m12_axi_arlen),
    .m_axi_rvalid(m12_axi_rvalid),
    .m_axi_rready(m12_axi_rready),
    .m_axi_rdata(m12_axi_rdata),
    .m_axi_rlast(m12_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid12),
    .m_axis_tready(rd_tready12),
    .m_axis_tlast(rd_tlast12),
    .m_axis_tdata(rd_tdata12)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_13
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[13]),
    .ctrl_addr_offset(in13),
    .ctrl_xfer_size_in_bytes(in_s13),
    .m_axi_arvalid(m13_axi_arvalid),
    .m_axi_arready(m13_axi_arready),
    .m_axi_araddr(m13_axi_araddr),
    .m_axi_arlen(m13_axi_arlen),
    .m_axi_rvalid(m13_axi_rvalid),
    .m_axi_rready(m13_axi_rready),
    .m_axi_rdata(m13_axi_rdata),
    .m_axi_rlast(m13_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid13),
    .m_axis_tready(rd_tready13),
    .m_axis_tlast(rd_tlast13),
    .m_axis_tdata(rd_tdata13)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_14
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[14]),
    .ctrl_addr_offset(in14),
    .ctrl_xfer_size_in_bytes(in_s14),
    .m_axi_arvalid(m14_axi_arvalid),
    .m_axi_arready(m14_axi_arready),
    .m_axi_araddr(m14_axi_araddr),
    .m_axi_arlen(m14_axi_arlen),
    .m_axi_rvalid(m14_axi_rvalid),
    .m_axi_rready(m14_axi_rready),
    .m_axi_rdata(m14_axi_rdata),
    .m_axi_rlast(m14_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid14),
    .m_axis_tready(rd_tready14),
    .m_axis_tlast(rd_tlast14),
    .m_axis_tdata(rd_tdata14)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_15
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[15]),
    .ctrl_addr_offset(in15),
    .ctrl_xfer_size_in_bytes(in_s15),
    .m_axi_arvalid(m15_axi_arvalid),
    .m_axi_arready(m15_axi_arready),
    .m_axi_araddr(m15_axi_araddr),
    .m_axi_arlen(m15_axi_arlen),
    .m_axi_rvalid(m15_axi_rvalid),
    .m_axi_rready(m15_axi_rready),
    .m_axi_rdata(m15_axi_rdata),
    .m_axi_rlast(m15_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid15),
    .m_axis_tready(rd_tready15),
    .m_axis_tlast(rd_tlast15),
    .m_axis_tdata(rd_tdata15)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_16
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[16]),
    .ctrl_addr_offset(in16),
    .ctrl_xfer_size_in_bytes(in_s16),
    .m_axi_arvalid(m16_axi_arvalid),
    .m_axi_arready(m16_axi_arready),
    .m_axi_araddr(m16_axi_araddr),
    .m_axi_arlen(m16_axi_arlen),
    .m_axi_rvalid(m16_axi_rvalid),
    .m_axi_rready(m16_axi_rready),
    .m_axi_rdata(m16_axi_rdata),
    .m_axi_rlast(m16_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid16),
    .m_axis_tready(rd_tready16),
    .m_axis_tlast(rd_tlast16),
    .m_axis_tdata(rd_tdata16)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_17
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[17]),
    .ctrl_addr_offset(in17),
    .ctrl_xfer_size_in_bytes(in_s17),
    .m_axi_arvalid(m17_axi_arvalid),
    .m_axi_arready(m17_axi_arready),
    .m_axi_araddr(m17_axi_araddr),
    .m_axi_arlen(m17_axi_arlen),
    .m_axi_rvalid(m17_axi_rvalid),
    .m_axi_rready(m17_axi_rready),
    .m_axi_rdata(m17_axi_rdata),
    .m_axi_rlast(m17_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid17),
    .m_axis_tready(rd_tready17),
    .m_axis_tlast(rd_tlast17),
    .m_axis_tdata(rd_tdata17)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_18
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[18]),
    .ctrl_addr_offset(in18),
    .ctrl_xfer_size_in_bytes(in_s18),
    .m_axi_arvalid(m18_axi_arvalid),
    .m_axi_arready(m18_axi_arready),
    .m_axi_araddr(m18_axi_araddr),
    .m_axi_arlen(m18_axi_arlen),
    .m_axi_rvalid(m18_axi_rvalid),
    .m_axi_rready(m18_axi_rready),
    .m_axi_rdata(m18_axi_rdata),
    .m_axi_rlast(m18_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid18),
    .m_axis_tready(rd_tready18),
    .m_axis_tlast(rd_tlast18),
    .m_axis_tdata(rd_tdata18)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_19
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[19]),
    .ctrl_addr_offset(in19),
    .ctrl_xfer_size_in_bytes(in_s19),
    .m_axi_arvalid(m19_axi_arvalid),
    .m_axi_arready(m19_axi_arready),
    .m_axi_araddr(m19_axi_araddr),
    .m_axi_arlen(m19_axi_arlen),
    .m_axi_rvalid(m19_axi_rvalid),
    .m_axi_rready(m19_axi_rready),
    .m_axi_rdata(m19_axi_rdata),
    .m_axi_rlast(m19_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid19),
    .m_axis_tready(rd_tready19),
    .m_axis_tlast(rd_tlast19),
    .m_axis_tdata(rd_tdata19)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_20
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[20]),
    .ctrl_addr_offset(in20),
    .ctrl_xfer_size_in_bytes(in_s20),
    .m_axi_arvalid(m20_axi_arvalid),
    .m_axi_arready(m20_axi_arready),
    .m_axi_araddr(m20_axi_araddr),
    .m_axi_arlen(m20_axi_arlen),
    .m_axi_rvalid(m20_axi_rvalid),
    .m_axi_rready(m20_axi_rready),
    .m_axi_rdata(m20_axi_rdata),
    .m_axi_rlast(m20_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid20),
    .m_axis_tready(rd_tready20),
    .m_axis_tlast(rd_tlast20),
    .m_axis_tdata(rd_tdata20)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_21
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[21]),
    .ctrl_addr_offset(in21),
    .ctrl_xfer_size_in_bytes(in_s21),
    .m_axi_arvalid(m21_axi_arvalid),
    .m_axi_arready(m21_axi_arready),
    .m_axi_araddr(m21_axi_araddr),
    .m_axi_arlen(m21_axi_arlen),
    .m_axi_rvalid(m21_axi_rvalid),
    .m_axi_rready(m21_axi_rready),
    .m_axi_rdata(m21_axi_rdata),
    .m_axi_rlast(m21_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid21),
    .m_axis_tready(rd_tready21),
    .m_axis_tlast(rd_tlast21),
    .m_axis_tdata(rd_tdata21)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_22
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[22]),
    .ctrl_addr_offset(in22),
    .ctrl_xfer_size_in_bytes(in_s22),
    .m_axi_arvalid(m22_axi_arvalid),
    .m_axi_arready(m22_axi_arready),
    .m_axi_araddr(m22_axi_araddr),
    .m_axi_arlen(m22_axi_arlen),
    .m_axi_rvalid(m22_axi_rvalid),
    .m_axi_rready(m22_axi_rready),
    .m_axi_rdata(m22_axi_rdata),
    .m_axi_rlast(m22_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid22),
    .m_axis_tready(rd_tready22),
    .m_axis_tlast(rd_tlast22),
    .m_axis_tdata(rd_tdata22)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_23
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[23]),
    .ctrl_addr_offset(in23),
    .ctrl_xfer_size_in_bytes(in_s23),
    .m_axi_arvalid(m23_axi_arvalid),
    .m_axi_arready(m23_axi_arready),
    .m_axi_araddr(m23_axi_araddr),
    .m_axi_arlen(m23_axi_arlen),
    .m_axi_rvalid(m23_axi_rvalid),
    .m_axi_rready(m23_axi_rready),
    .m_axi_rdata(m23_axi_rdata),
    .m_axi_rlast(m23_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid23),
    .m_axis_tready(rd_tready23),
    .m_axis_tlast(rd_tlast23),
    .m_axis_tdata(rd_tdata23)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_24
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[24]),
    .ctrl_addr_offset(in24),
    .ctrl_xfer_size_in_bytes(in_s24),
    .m_axi_arvalid(m24_axi_arvalid),
    .m_axi_arready(m24_axi_arready),
    .m_axi_araddr(m24_axi_araddr),
    .m_axi_arlen(m24_axi_arlen),
    .m_axi_rvalid(m24_axi_rvalid),
    .m_axi_rready(m24_axi_rready),
    .m_axi_rdata(m24_axi_rdata),
    .m_axi_rlast(m24_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid24),
    .m_axis_tready(rd_tready24),
    .m_axis_tlast(rd_tlast24),
    .m_axis_tdata(rd_tdata24)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_25
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[25]),
    .ctrl_addr_offset(in25),
    .ctrl_xfer_size_in_bytes(in_s25),
    .m_axi_arvalid(m25_axi_arvalid),
    .m_axi_arready(m25_axi_arready),
    .m_axi_araddr(m25_axi_araddr),
    .m_axi_arlen(m25_axi_arlen),
    .m_axi_rvalid(m25_axi_rvalid),
    .m_axi_rready(m25_axi_rready),
    .m_axi_rdata(m25_axi_rdata),
    .m_axi_rlast(m25_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid25),
    .m_axis_tready(rd_tready25),
    .m_axis_tlast(rd_tlast25),
    .m_axis_tdata(rd_tdata25)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_26
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[26]),
    .ctrl_addr_offset(in26),
    .ctrl_xfer_size_in_bytes(in_s26),
    .m_axi_arvalid(m26_axi_arvalid),
    .m_axi_arready(m26_axi_arready),
    .m_axi_araddr(m26_axi_araddr),
    .m_axi_arlen(m26_axi_arlen),
    .m_axi_rvalid(m26_axi_rvalid),
    .m_axi_rready(m26_axi_rready),
    .m_axi_rdata(m26_axi_rdata),
    .m_axi_rlast(m26_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid26),
    .m_axis_tready(rd_tready26),
    .m_axis_tlast(rd_tlast26),
    .m_axis_tdata(rd_tdata26)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_27
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[27]),
    .ctrl_addr_offset(in27),
    .ctrl_xfer_size_in_bytes(in_s27),
    .m_axi_arvalid(m27_axi_arvalid),
    .m_axi_arready(m27_axi_arready),
    .m_axi_araddr(m27_axi_araddr),
    .m_axi_arlen(m27_axi_arlen),
    .m_axi_rvalid(m27_axi_rvalid),
    .m_axi_rready(m27_axi_rready),
    .m_axi_rdata(m27_axi_rdata),
    .m_axi_rlast(m27_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid27),
    .m_axis_tready(rd_tready27),
    .m_axis_tlast(rd_tlast27),
    .m_axis_tdata(rd_tdata27)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_28
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[28]),
    .ctrl_addr_offset(in28),
    .ctrl_xfer_size_in_bytes(in_s28),
    .m_axi_arvalid(m28_axi_arvalid),
    .m_axi_arready(m28_axi_arready),
    .m_axi_araddr(m28_axi_araddr),
    .m_axi_arlen(m28_axi_arlen),
    .m_axi_rvalid(m28_axi_rvalid),
    .m_axi_rready(m28_axi_rready),
    .m_axi_rdata(m28_axi_rdata),
    .m_axi_rlast(m28_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid28),
    .m_axis_tready(rd_tready28),
    .m_axis_tlast(rd_tlast28),
    .m_axis_tdata(rd_tdata28)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_29
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[29]),
    .ctrl_addr_offset(in29),
    .ctrl_xfer_size_in_bytes(in_s29),
    .m_axi_arvalid(m29_axi_arvalid),
    .m_axi_arready(m29_axi_arready),
    .m_axi_araddr(m29_axi_araddr),
    .m_axi_arlen(m29_axi_arlen),
    .m_axi_rvalid(m29_axi_rvalid),
    .m_axi_rready(m29_axi_rready),
    .m_axi_rdata(m29_axi_rdata),
    .m_axi_rlast(m29_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid29),
    .m_axis_tready(rd_tready29),
    .m_axis_tlast(rd_tlast29),
    .m_axis_tdata(rd_tdata29)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_30
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[30]),
    .ctrl_addr_offset(in30),
    .ctrl_xfer_size_in_bytes(in_s30),
    .m_axi_arvalid(m30_axi_arvalid),
    .m_axi_arready(m30_axi_arready),
    .m_axi_araddr(m30_axi_araddr),
    .m_axi_arlen(m30_axi_arlen),
    .m_axi_rvalid(m30_axi_rvalid),
    .m_axi_rready(m30_axi_rready),
    .m_axi_rdata(m30_axi_rdata),
    .m_axi_rlast(m30_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid30),
    .m_axis_tready(rd_tready30),
    .m_axis_tlast(rd_tlast30),
    .m_axis_tdata(rd_tdata30)
  );


  axi_reader_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_RD_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_reader_31
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(rd_ctrl_done[31]),
    .ctrl_addr_offset(in31),
    .ctrl_xfer_size_in_bytes(in_s31),
    .m_axi_arvalid(m31_axi_arvalid),
    .m_axi_arready(m31_axi_arready),
    .m_axi_araddr(m31_axi_araddr),
    .m_axi_arlen(m31_axi_arlen),
    .m_axi_rvalid(m31_axi_rvalid),
    .m_axi_rready(m31_axi_rready),
    .m_axi_rdata(m31_axi_rdata),
    .m_axi_rlast(m31_axi_rlast),
    .m_axis_aclk(ap_clk),
    .m_axis_areset(areset),
    .m_axis_tvalid(rd_tvalid31),
    .m_axis_tready(rd_tready31),
    .m_axis_tlast(rd_tlast31),
    .m_axis_tdata(rd_tdata31)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_0
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[0]),
    .ctrl_addr_offset(out0),
    .ctrl_xfer_size_in_bytes(out_s0),
    .m_axi_awvalid(m00_axi_awvalid),
    .m_axi_awready(m00_axi_awready),
    .m_axi_awaddr(m00_axi_awaddr),
    .m_axi_awlen(m00_axi_awlen),
    .m_axi_wvalid(m00_axi_wvalid),
    .m_axi_wready(m00_axi_wready),
    .m_axi_wdata(m00_axi_wdata),
    .m_axi_wstrb(m00_axi_wstrb),
    .m_axi_wlast(m00_axi_wlast),
    .m_axi_bvalid(m00_axi_bvalid),
    .m_axi_bready(m00_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid0),
    .s_axis_tready(wr_tready0),
    .s_axis_tdata(wr_tdata0)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_1
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[1]),
    .ctrl_addr_offset(out1),
    .ctrl_xfer_size_in_bytes(out_s1),
    .m_axi_awvalid(m01_axi_awvalid),
    .m_axi_awready(m01_axi_awready),
    .m_axi_awaddr(m01_axi_awaddr),
    .m_axi_awlen(m01_axi_awlen),
    .m_axi_wvalid(m01_axi_wvalid),
    .m_axi_wready(m01_axi_wready),
    .m_axi_wdata(m01_axi_wdata),
    .m_axi_wstrb(m01_axi_wstrb),
    .m_axi_wlast(m01_axi_wlast),
    .m_axi_bvalid(m01_axi_bvalid),
    .m_axi_bready(m01_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid1),
    .s_axis_tready(wr_tready1),
    .s_axis_tdata(wr_tdata1)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_2
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[2]),
    .ctrl_addr_offset(out2),
    .ctrl_xfer_size_in_bytes(out_s2),
    .m_axi_awvalid(m02_axi_awvalid),
    .m_axi_awready(m02_axi_awready),
    .m_axi_awaddr(m02_axi_awaddr),
    .m_axi_awlen(m02_axi_awlen),
    .m_axi_wvalid(m02_axi_wvalid),
    .m_axi_wready(m02_axi_wready),
    .m_axi_wdata(m02_axi_wdata),
    .m_axi_wstrb(m02_axi_wstrb),
    .m_axi_wlast(m02_axi_wlast),
    .m_axi_bvalid(m02_axi_bvalid),
    .m_axi_bready(m02_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid2),
    .s_axis_tready(wr_tready2),
    .s_axis_tdata(wr_tdata2)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_3
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[3]),
    .ctrl_addr_offset(out3),
    .ctrl_xfer_size_in_bytes(out_s3),
    .m_axi_awvalid(m03_axi_awvalid),
    .m_axi_awready(m03_axi_awready),
    .m_axi_awaddr(m03_axi_awaddr),
    .m_axi_awlen(m03_axi_awlen),
    .m_axi_wvalid(m03_axi_wvalid),
    .m_axi_wready(m03_axi_wready),
    .m_axi_wdata(m03_axi_wdata),
    .m_axi_wstrb(m03_axi_wstrb),
    .m_axi_wlast(m03_axi_wlast),
    .m_axi_bvalid(m03_axi_bvalid),
    .m_axi_bready(m03_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid3),
    .s_axis_tready(wr_tready3),
    .s_axis_tdata(wr_tdata3)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_4
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[4]),
    .ctrl_addr_offset(out4),
    .ctrl_xfer_size_in_bytes(out_s4),
    .m_axi_awvalid(m04_axi_awvalid),
    .m_axi_awready(m04_axi_awready),
    .m_axi_awaddr(m04_axi_awaddr),
    .m_axi_awlen(m04_axi_awlen),
    .m_axi_wvalid(m04_axi_wvalid),
    .m_axi_wready(m04_axi_wready),
    .m_axi_wdata(m04_axi_wdata),
    .m_axi_wstrb(m04_axi_wstrb),
    .m_axi_wlast(m04_axi_wlast),
    .m_axi_bvalid(m04_axi_bvalid),
    .m_axi_bready(m04_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid4),
    .s_axis_tready(wr_tready4),
    .s_axis_tdata(wr_tdata4)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_5
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[5]),
    .ctrl_addr_offset(out5),
    .ctrl_xfer_size_in_bytes(out_s5),
    .m_axi_awvalid(m05_axi_awvalid),
    .m_axi_awready(m05_axi_awready),
    .m_axi_awaddr(m05_axi_awaddr),
    .m_axi_awlen(m05_axi_awlen),
    .m_axi_wvalid(m05_axi_wvalid),
    .m_axi_wready(m05_axi_wready),
    .m_axi_wdata(m05_axi_wdata),
    .m_axi_wstrb(m05_axi_wstrb),
    .m_axi_wlast(m05_axi_wlast),
    .m_axi_bvalid(m05_axi_bvalid),
    .m_axi_bready(m05_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid5),
    .s_axis_tready(wr_tready5),
    .s_axis_tdata(wr_tdata5)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_6
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[6]),
    .ctrl_addr_offset(out6),
    .ctrl_xfer_size_in_bytes(out_s6),
    .m_axi_awvalid(m06_axi_awvalid),
    .m_axi_awready(m06_axi_awready),
    .m_axi_awaddr(m06_axi_awaddr),
    .m_axi_awlen(m06_axi_awlen),
    .m_axi_wvalid(m06_axi_wvalid),
    .m_axi_wready(m06_axi_wready),
    .m_axi_wdata(m06_axi_wdata),
    .m_axi_wstrb(m06_axi_wstrb),
    .m_axi_wlast(m06_axi_wlast),
    .m_axi_bvalid(m06_axi_bvalid),
    .m_axi_bready(m06_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid6),
    .s_axis_tready(wr_tready6),
    .s_axis_tdata(wr_tdata6)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_7
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[7]),
    .ctrl_addr_offset(out7),
    .ctrl_xfer_size_in_bytes(out_s7),
    .m_axi_awvalid(m07_axi_awvalid),
    .m_axi_awready(m07_axi_awready),
    .m_axi_awaddr(m07_axi_awaddr),
    .m_axi_awlen(m07_axi_awlen),
    .m_axi_wvalid(m07_axi_wvalid),
    .m_axi_wready(m07_axi_wready),
    .m_axi_wdata(m07_axi_wdata),
    .m_axi_wstrb(m07_axi_wstrb),
    .m_axi_wlast(m07_axi_wlast),
    .m_axi_bvalid(m07_axi_bvalid),
    .m_axi_bready(m07_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid7),
    .s_axis_tready(wr_tready7),
    .s_axis_tdata(wr_tdata7)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_8
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[8]),
    .ctrl_addr_offset(out8),
    .ctrl_xfer_size_in_bytes(out_s8),
    .m_axi_awvalid(m08_axi_awvalid),
    .m_axi_awready(m08_axi_awready),
    .m_axi_awaddr(m08_axi_awaddr),
    .m_axi_awlen(m08_axi_awlen),
    .m_axi_wvalid(m08_axi_wvalid),
    .m_axi_wready(m08_axi_wready),
    .m_axi_wdata(m08_axi_wdata),
    .m_axi_wstrb(m08_axi_wstrb),
    .m_axi_wlast(m08_axi_wlast),
    .m_axi_bvalid(m08_axi_bvalid),
    .m_axi_bready(m08_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid8),
    .s_axis_tready(wr_tready8),
    .s_axis_tdata(wr_tdata8)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_9
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[9]),
    .ctrl_addr_offset(out9),
    .ctrl_xfer_size_in_bytes(out_s9),
    .m_axi_awvalid(m09_axi_awvalid),
    .m_axi_awready(m09_axi_awready),
    .m_axi_awaddr(m09_axi_awaddr),
    .m_axi_awlen(m09_axi_awlen),
    .m_axi_wvalid(m09_axi_wvalid),
    .m_axi_wready(m09_axi_wready),
    .m_axi_wdata(m09_axi_wdata),
    .m_axi_wstrb(m09_axi_wstrb),
    .m_axi_wlast(m09_axi_wlast),
    .m_axi_bvalid(m09_axi_bvalid),
    .m_axi_bready(m09_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid9),
    .s_axis_tready(wr_tready9),
    .s_axis_tdata(wr_tdata9)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_10
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[10]),
    .ctrl_addr_offset(out10),
    .ctrl_xfer_size_in_bytes(out_s10),
    .m_axi_awvalid(m10_axi_awvalid),
    .m_axi_awready(m10_axi_awready),
    .m_axi_awaddr(m10_axi_awaddr),
    .m_axi_awlen(m10_axi_awlen),
    .m_axi_wvalid(m10_axi_wvalid),
    .m_axi_wready(m10_axi_wready),
    .m_axi_wdata(m10_axi_wdata),
    .m_axi_wstrb(m10_axi_wstrb),
    .m_axi_wlast(m10_axi_wlast),
    .m_axi_bvalid(m10_axi_bvalid),
    .m_axi_bready(m10_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid10),
    .s_axis_tready(wr_tready10),
    .s_axis_tdata(wr_tdata10)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_11
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[11]),
    .ctrl_addr_offset(out11),
    .ctrl_xfer_size_in_bytes(out_s11),
    .m_axi_awvalid(m11_axi_awvalid),
    .m_axi_awready(m11_axi_awready),
    .m_axi_awaddr(m11_axi_awaddr),
    .m_axi_awlen(m11_axi_awlen),
    .m_axi_wvalid(m11_axi_wvalid),
    .m_axi_wready(m11_axi_wready),
    .m_axi_wdata(m11_axi_wdata),
    .m_axi_wstrb(m11_axi_wstrb),
    .m_axi_wlast(m11_axi_wlast),
    .m_axi_bvalid(m11_axi_bvalid),
    .m_axi_bready(m11_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid11),
    .s_axis_tready(wr_tready11),
    .s_axis_tdata(wr_tdata11)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_12
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[12]),
    .ctrl_addr_offset(out12),
    .ctrl_xfer_size_in_bytes(out_s12),
    .m_axi_awvalid(m12_axi_awvalid),
    .m_axi_awready(m12_axi_awready),
    .m_axi_awaddr(m12_axi_awaddr),
    .m_axi_awlen(m12_axi_awlen),
    .m_axi_wvalid(m12_axi_wvalid),
    .m_axi_wready(m12_axi_wready),
    .m_axi_wdata(m12_axi_wdata),
    .m_axi_wstrb(m12_axi_wstrb),
    .m_axi_wlast(m12_axi_wlast),
    .m_axi_bvalid(m12_axi_bvalid),
    .m_axi_bready(m12_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid12),
    .s_axis_tready(wr_tready12),
    .s_axis_tdata(wr_tdata12)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_13
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[13]),
    .ctrl_addr_offset(out13),
    .ctrl_xfer_size_in_bytes(out_s13),
    .m_axi_awvalid(m13_axi_awvalid),
    .m_axi_awready(m13_axi_awready),
    .m_axi_awaddr(m13_axi_awaddr),
    .m_axi_awlen(m13_axi_awlen),
    .m_axi_wvalid(m13_axi_wvalid),
    .m_axi_wready(m13_axi_wready),
    .m_axi_wdata(m13_axi_wdata),
    .m_axi_wstrb(m13_axi_wstrb),
    .m_axi_wlast(m13_axi_wlast),
    .m_axi_bvalid(m13_axi_bvalid),
    .m_axi_bready(m13_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid13),
    .s_axis_tready(wr_tready13),
    .s_axis_tdata(wr_tdata13)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_14
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[14]),
    .ctrl_addr_offset(out14),
    .ctrl_xfer_size_in_bytes(out_s14),
    .m_axi_awvalid(m14_axi_awvalid),
    .m_axi_awready(m14_axi_awready),
    .m_axi_awaddr(m14_axi_awaddr),
    .m_axi_awlen(m14_axi_awlen),
    .m_axi_wvalid(m14_axi_wvalid),
    .m_axi_wready(m14_axi_wready),
    .m_axi_wdata(m14_axi_wdata),
    .m_axi_wstrb(m14_axi_wstrb),
    .m_axi_wlast(m14_axi_wlast),
    .m_axi_bvalid(m14_axi_bvalid),
    .m_axi_bready(m14_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid14),
    .s_axis_tready(wr_tready14),
    .s_axis_tdata(wr_tdata14)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_15
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[15]),
    .ctrl_addr_offset(out15),
    .ctrl_xfer_size_in_bytes(out_s15),
    .m_axi_awvalid(m15_axi_awvalid),
    .m_axi_awready(m15_axi_awready),
    .m_axi_awaddr(m15_axi_awaddr),
    .m_axi_awlen(m15_axi_awlen),
    .m_axi_wvalid(m15_axi_wvalid),
    .m_axi_wready(m15_axi_wready),
    .m_axi_wdata(m15_axi_wdata),
    .m_axi_wstrb(m15_axi_wstrb),
    .m_axi_wlast(m15_axi_wlast),
    .m_axi_bvalid(m15_axi_bvalid),
    .m_axi_bready(m15_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid15),
    .s_axis_tready(wr_tready15),
    .s_axis_tdata(wr_tdata15)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_16
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[16]),
    .ctrl_addr_offset(out16),
    .ctrl_xfer_size_in_bytes(out_s16),
    .m_axi_awvalid(m16_axi_awvalid),
    .m_axi_awready(m16_axi_awready),
    .m_axi_awaddr(m16_axi_awaddr),
    .m_axi_awlen(m16_axi_awlen),
    .m_axi_wvalid(m16_axi_wvalid),
    .m_axi_wready(m16_axi_wready),
    .m_axi_wdata(m16_axi_wdata),
    .m_axi_wstrb(m16_axi_wstrb),
    .m_axi_wlast(m16_axi_wlast),
    .m_axi_bvalid(m16_axi_bvalid),
    .m_axi_bready(m16_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid16),
    .s_axis_tready(wr_tready16),
    .s_axis_tdata(wr_tdata16)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_17
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[17]),
    .ctrl_addr_offset(out17),
    .ctrl_xfer_size_in_bytes(out_s17),
    .m_axi_awvalid(m17_axi_awvalid),
    .m_axi_awready(m17_axi_awready),
    .m_axi_awaddr(m17_axi_awaddr),
    .m_axi_awlen(m17_axi_awlen),
    .m_axi_wvalid(m17_axi_wvalid),
    .m_axi_wready(m17_axi_wready),
    .m_axi_wdata(m17_axi_wdata),
    .m_axi_wstrb(m17_axi_wstrb),
    .m_axi_wlast(m17_axi_wlast),
    .m_axi_bvalid(m17_axi_bvalid),
    .m_axi_bready(m17_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid17),
    .s_axis_tready(wr_tready17),
    .s_axis_tdata(wr_tdata17)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_18
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[18]),
    .ctrl_addr_offset(out18),
    .ctrl_xfer_size_in_bytes(out_s18),
    .m_axi_awvalid(m18_axi_awvalid),
    .m_axi_awready(m18_axi_awready),
    .m_axi_awaddr(m18_axi_awaddr),
    .m_axi_awlen(m18_axi_awlen),
    .m_axi_wvalid(m18_axi_wvalid),
    .m_axi_wready(m18_axi_wready),
    .m_axi_wdata(m18_axi_wdata),
    .m_axi_wstrb(m18_axi_wstrb),
    .m_axi_wlast(m18_axi_wlast),
    .m_axi_bvalid(m18_axi_bvalid),
    .m_axi_bready(m18_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid18),
    .s_axis_tready(wr_tready18),
    .s_axis_tdata(wr_tdata18)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_19
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[19]),
    .ctrl_addr_offset(out19),
    .ctrl_xfer_size_in_bytes(out_s19),
    .m_axi_awvalid(m19_axi_awvalid),
    .m_axi_awready(m19_axi_awready),
    .m_axi_awaddr(m19_axi_awaddr),
    .m_axi_awlen(m19_axi_awlen),
    .m_axi_wvalid(m19_axi_wvalid),
    .m_axi_wready(m19_axi_wready),
    .m_axi_wdata(m19_axi_wdata),
    .m_axi_wstrb(m19_axi_wstrb),
    .m_axi_wlast(m19_axi_wlast),
    .m_axi_bvalid(m19_axi_bvalid),
    .m_axi_bready(m19_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid19),
    .s_axis_tready(wr_tready19),
    .s_axis_tdata(wr_tdata19)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_20
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[20]),
    .ctrl_addr_offset(out20),
    .ctrl_xfer_size_in_bytes(out_s20),
    .m_axi_awvalid(m20_axi_awvalid),
    .m_axi_awready(m20_axi_awready),
    .m_axi_awaddr(m20_axi_awaddr),
    .m_axi_awlen(m20_axi_awlen),
    .m_axi_wvalid(m20_axi_wvalid),
    .m_axi_wready(m20_axi_wready),
    .m_axi_wdata(m20_axi_wdata),
    .m_axi_wstrb(m20_axi_wstrb),
    .m_axi_wlast(m20_axi_wlast),
    .m_axi_bvalid(m20_axi_bvalid),
    .m_axi_bready(m20_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid20),
    .s_axis_tready(wr_tready20),
    .s_axis_tdata(wr_tdata20)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_21
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[21]),
    .ctrl_addr_offset(out21),
    .ctrl_xfer_size_in_bytes(out_s21),
    .m_axi_awvalid(m21_axi_awvalid),
    .m_axi_awready(m21_axi_awready),
    .m_axi_awaddr(m21_axi_awaddr),
    .m_axi_awlen(m21_axi_awlen),
    .m_axi_wvalid(m21_axi_wvalid),
    .m_axi_wready(m21_axi_wready),
    .m_axi_wdata(m21_axi_wdata),
    .m_axi_wstrb(m21_axi_wstrb),
    .m_axi_wlast(m21_axi_wlast),
    .m_axi_bvalid(m21_axi_bvalid),
    .m_axi_bready(m21_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid21),
    .s_axis_tready(wr_tready21),
    .s_axis_tdata(wr_tdata21)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_22
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[22]),
    .ctrl_addr_offset(out22),
    .ctrl_xfer_size_in_bytes(out_s22),
    .m_axi_awvalid(m22_axi_awvalid),
    .m_axi_awready(m22_axi_awready),
    .m_axi_awaddr(m22_axi_awaddr),
    .m_axi_awlen(m22_axi_awlen),
    .m_axi_wvalid(m22_axi_wvalid),
    .m_axi_wready(m22_axi_wready),
    .m_axi_wdata(m22_axi_wdata),
    .m_axi_wstrb(m22_axi_wstrb),
    .m_axi_wlast(m22_axi_wlast),
    .m_axi_bvalid(m22_axi_bvalid),
    .m_axi_bready(m22_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid22),
    .s_axis_tready(wr_tready22),
    .s_axis_tdata(wr_tdata22)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_23
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[23]),
    .ctrl_addr_offset(out23),
    .ctrl_xfer_size_in_bytes(out_s23),
    .m_axi_awvalid(m23_axi_awvalid),
    .m_axi_awready(m23_axi_awready),
    .m_axi_awaddr(m23_axi_awaddr),
    .m_axi_awlen(m23_axi_awlen),
    .m_axi_wvalid(m23_axi_wvalid),
    .m_axi_wready(m23_axi_wready),
    .m_axi_wdata(m23_axi_wdata),
    .m_axi_wstrb(m23_axi_wstrb),
    .m_axi_wlast(m23_axi_wlast),
    .m_axi_bvalid(m23_axi_bvalid),
    .m_axi_bready(m23_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid23),
    .s_axis_tready(wr_tready23),
    .s_axis_tdata(wr_tdata23)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_24
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[24]),
    .ctrl_addr_offset(out24),
    .ctrl_xfer_size_in_bytes(out_s24),
    .m_axi_awvalid(m24_axi_awvalid),
    .m_axi_awready(m24_axi_awready),
    .m_axi_awaddr(m24_axi_awaddr),
    .m_axi_awlen(m24_axi_awlen),
    .m_axi_wvalid(m24_axi_wvalid),
    .m_axi_wready(m24_axi_wready),
    .m_axi_wdata(m24_axi_wdata),
    .m_axi_wstrb(m24_axi_wstrb),
    .m_axi_wlast(m24_axi_wlast),
    .m_axi_bvalid(m24_axi_bvalid),
    .m_axi_bready(m24_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid24),
    .s_axis_tready(wr_tready24),
    .s_axis_tdata(wr_tdata24)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_25
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[25]),
    .ctrl_addr_offset(out25),
    .ctrl_xfer_size_in_bytes(out_s25),
    .m_axi_awvalid(m25_axi_awvalid),
    .m_axi_awready(m25_axi_awready),
    .m_axi_awaddr(m25_axi_awaddr),
    .m_axi_awlen(m25_axi_awlen),
    .m_axi_wvalid(m25_axi_wvalid),
    .m_axi_wready(m25_axi_wready),
    .m_axi_wdata(m25_axi_wdata),
    .m_axi_wstrb(m25_axi_wstrb),
    .m_axi_wlast(m25_axi_wlast),
    .m_axi_bvalid(m25_axi_bvalid),
    .m_axi_bready(m25_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid25),
    .s_axis_tready(wr_tready25),
    .s_axis_tdata(wr_tdata25)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_26
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[26]),
    .ctrl_addr_offset(out26),
    .ctrl_xfer_size_in_bytes(out_s26),
    .m_axi_awvalid(m26_axi_awvalid),
    .m_axi_awready(m26_axi_awready),
    .m_axi_awaddr(m26_axi_awaddr),
    .m_axi_awlen(m26_axi_awlen),
    .m_axi_wvalid(m26_axi_wvalid),
    .m_axi_wready(m26_axi_wready),
    .m_axi_wdata(m26_axi_wdata),
    .m_axi_wstrb(m26_axi_wstrb),
    .m_axi_wlast(m26_axi_wlast),
    .m_axi_bvalid(m26_axi_bvalid),
    .m_axi_bready(m26_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid26),
    .s_axis_tready(wr_tready26),
    .s_axis_tdata(wr_tdata26)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_27
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[27]),
    .ctrl_addr_offset(out27),
    .ctrl_xfer_size_in_bytes(out_s27),
    .m_axi_awvalid(m27_axi_awvalid),
    .m_axi_awready(m27_axi_awready),
    .m_axi_awaddr(m27_axi_awaddr),
    .m_axi_awlen(m27_axi_awlen),
    .m_axi_wvalid(m27_axi_wvalid),
    .m_axi_wready(m27_axi_wready),
    .m_axi_wdata(m27_axi_wdata),
    .m_axi_wstrb(m27_axi_wstrb),
    .m_axi_wlast(m27_axi_wlast),
    .m_axi_bvalid(m27_axi_bvalid),
    .m_axi_bready(m27_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid27),
    .s_axis_tready(wr_tready27),
    .s_axis_tdata(wr_tdata27)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_28
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[28]),
    .ctrl_addr_offset(out28),
    .ctrl_xfer_size_in_bytes(out_s28),
    .m_axi_awvalid(m28_axi_awvalid),
    .m_axi_awready(m28_axi_awready),
    .m_axi_awaddr(m28_axi_awaddr),
    .m_axi_awlen(m28_axi_awlen),
    .m_axi_wvalid(m28_axi_wvalid),
    .m_axi_wready(m28_axi_wready),
    .m_axi_wdata(m28_axi_wdata),
    .m_axi_wstrb(m28_axi_wstrb),
    .m_axi_wlast(m28_axi_wlast),
    .m_axi_bvalid(m28_axi_bvalid),
    .m_axi_bready(m28_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid28),
    .s_axis_tready(wr_tready28),
    .s_axis_tdata(wr_tdata28)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_29
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[29]),
    .ctrl_addr_offset(out29),
    .ctrl_xfer_size_in_bytes(out_s29),
    .m_axi_awvalid(m29_axi_awvalid),
    .m_axi_awready(m29_axi_awready),
    .m_axi_awaddr(m29_axi_awaddr),
    .m_axi_awlen(m29_axi_awlen),
    .m_axi_wvalid(m29_axi_wvalid),
    .m_axi_wready(m29_axi_wready),
    .m_axi_wdata(m29_axi_wdata),
    .m_axi_wstrb(m29_axi_wstrb),
    .m_axi_wlast(m29_axi_wlast),
    .m_axi_bvalid(m29_axi_bvalid),
    .m_axi_bready(m29_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid29),
    .s_axis_tready(wr_tready29),
    .s_axis_tdata(wr_tdata29)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_30
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[30]),
    .ctrl_addr_offset(out30),
    .ctrl_xfer_size_in_bytes(out_s30),
    .m_axi_awvalid(m30_axi_awvalid),
    .m_axi_awready(m30_axi_awready),
    .m_axi_awaddr(m30_axi_awaddr),
    .m_axi_awlen(m30_axi_awlen),
    .m_axi_wvalid(m30_axi_wvalid),
    .m_axi_wready(m30_axi_wready),
    .m_axi_wdata(m30_axi_wdata),
    .m_axi_wstrb(m30_axi_wstrb),
    .m_axi_wlast(m30_axi_wlast),
    .m_axi_bvalid(m30_axi_bvalid),
    .m_axi_bready(m30_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid30),
    .s_axis_tready(wr_tready30),
    .s_axis_tdata(wr_tdata30)
  );


  axi_writer_wrapper
  #(
    .C_M_AXI_ADDR_WIDTH(C_M_AXI_ADDR_WIDTH),
    .C_M_AXI_DATA_WIDTH(C_M_AXI_DATA_WIDTH),
    .C_XFER_SIZE_WIDTH(32),
    .C_MAX_OUTSTANDING(LP_WR_MAX_OUTSTANDING),
    .C_INCLUDE_DATA_FIFO(1)
  )
  axi_writer_31
  (
    .aclk(ap_clk),
    .areset(areset),
    .ctrl_start(ap_start_pulse),
    .ctrl_done(wr_ctrl_done[31]),
    .ctrl_addr_offset(out31),
    .ctrl_xfer_size_in_bytes(out_s31),
    .m_axi_awvalid(m31_axi_awvalid),
    .m_axi_awready(m31_axi_awready),
    .m_axi_awaddr(m31_axi_awaddr),
    .m_axi_awlen(m31_axi_awlen),
    .m_axi_wvalid(m31_axi_wvalid),
    .m_axi_wready(m31_axi_wready),
    .m_axi_wdata(m31_axi_wdata),
    .m_axi_wstrb(m31_axi_wstrb),
    .m_axi_wlast(m31_axi_wlast),
    .m_axi_bvalid(m31_axi_bvalid),
    .m_axi_bready(m31_axi_bready),
    .s_axis_aclk(ap_clk),
    .s_axis_areset(areset),
    .s_axis_tvalid(wr_tvalid31),
    .s_axis_tready(wr_tready31),
    .s_axis_tdata(wr_tdata31)
  );


  m_accelerator
  acc
  (
    .clk(ap_clk),
    .rst(areset),
    .start(user_start),
    .acc_user_done_rd_data(acc_user_done_rd_data),
    .acc_user_done_wr_data(acc_user_done_wr_data),
    .acc_user_request_read(acc_user_request_read),
    .acc_user_read_data_valid(acc_user_read_data_valid),
    .acc_user_read_data(acc_user_read_data),
    .acc_user_available_write(acc_user_available_write),
    .acc_user_request_write(acc_user_request_write),
    .acc_user_write_data(acc_user_write_data),
    .acc_user_done(acc_user_done)
  );


  initial begin
    reset = 1'b1;
    ap_idle_r = 1'b1;
    ap_done_r = 0;
    acc_user_done_rd_data = 0;
    acc_user_done_wr_data = 0;
    fsm_reset = FSM_STATE_START;
    areset = 1'b1;
    ap_start_pulse = 0;
    user_start = 0;
  end


endmodule



module axi_reader_wrapper #
(
  parameter C_M_AXI_ADDR_WIDTH = 64,
  parameter C_M_AXI_DATA_WIDTH = 256,
  parameter C_XFER_SIZE_WIDTH = 64,
  parameter C_MAX_OUTSTANDING = 16,
  parameter C_INCLUDE_DATA_FIFO = 1
)
(
  input aclk,
  input areset,
  input ctrl_start,
  output ctrl_done,
  input [C_M_AXI_ADDR_WIDTH-1:0] ctrl_addr_offset,
  input [C_XFER_SIZE_WIDTH-1:0] ctrl_xfer_size_in_bytes,
  output m_axi_arvalid,
  input m_axi_arready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m_axi_araddr,
  output [8-1:0] m_axi_arlen,
  input m_axi_rvalid,
  output m_axi_rready,
  input [C_M_AXI_DATA_WIDTH-1:0] m_axi_rdata,
  input m_axi_rlast,
  input m_axis_aclk,
  input m_axis_areset,
  output m_axis_tvalid,
  input m_axis_tready,
  output [C_M_AXI_DATA_WIDTH-1:0] m_axis_tdata,
  output m_axis_tlast
);

  axi_reader #(
            .C_M_AXI_ADDR_WIDTH  ( C_M_AXI_ADDR_WIDTH  ) ,
            .C_M_AXI_DATA_WIDTH  ( C_M_AXI_DATA_WIDTH  ) ,
            .C_XFER_SIZE_WIDTH   ( C_XFER_SIZE_WIDTH   ) ,
            .C_MAX_OUTSTANDING   ( C_MAX_OUTSTANDING   ) ,
            .C_INCLUDE_DATA_FIFO ( C_INCLUDE_DATA_FIFO )
          )
          inst_axi_reader (
            .aclk                    ( aclk                   ) ,
            .areset                  ( areset                 ) ,
            .ctrl_start              ( ctrl_start             ) ,
            .ctrl_done               ( ctrl_done              ) ,
            .ctrl_addr_offset        ( ctrl_addr_offset       ) ,
            .ctrl_xfer_size_in_bytes ( ctrl_xfer_size_in_bytes) ,
            .m_axi_arvalid           ( m_axi_arvalid          ) ,
            .m_axi_arready           ( m_axi_arready          ) ,
            .m_axi_araddr            ( m_axi_araddr           ) ,
            .m_axi_arlen             ( m_axi_arlen            ) ,
            .m_axi_rvalid            ( m_axi_rvalid           ) ,
            .m_axi_rready            ( m_axi_rready           ) ,
            .m_axi_rdata             ( m_axi_rdata            ) ,
            .m_axi_rlast             ( m_axi_rlast            ) ,
            .m_axis_aclk             ( m_axis_aclk            ) ,
            .m_axis_areset           ( m_axis_areset          ) ,
            .m_axis_tvalid           ( m_axis_tvalid          ) ,
            .m_axis_tready           ( m_axis_tready          ) ,
            .m_axis_tlast            ( m_axis_tlast           ) ,
            .m_axis_tdata            ( m_axis_tdata           )
          );

endmodule



module axi_writer_wrapper #
(
  parameter C_M_AXI_ADDR_WIDTH = 64,
  parameter C_M_AXI_DATA_WIDTH = 256,
  parameter C_XFER_SIZE_WIDTH = 64,
  parameter C_MAX_OUTSTANDING = 16,
  parameter C_INCLUDE_DATA_FIFO = 1
)
(
  input aclk,
  input areset,
  input ctrl_start,
  output ctrl_done,
  input [C_M_AXI_ADDR_WIDTH-1:0] ctrl_addr_offset,
  input [C_XFER_SIZE_WIDTH-1:0] ctrl_xfer_size_in_bytes,
  output m_axi_awvalid,
  input m_axi_awready,
  output [C_M_AXI_ADDR_WIDTH-1:0] m_axi_awaddr,
  output [8-1:0] m_axi_awlen,
  output m_axi_wvalid,
  input m_axi_wready,
  output [C_M_AXI_DATA_WIDTH-1:0] m_axi_wdata,
  output [C_M_AXI_DATA_WIDTH/8-1:0] m_axi_wstrb,
  output m_axi_wlast,
  input m_axi_bvalid,
  output m_axi_bready,
  input s_axis_aclk,
  input s_axis_areset,
  input s_axis_tvalid,
  output s_axis_tready,
  input [C_M_AXI_DATA_WIDTH-1:0] s_axis_tdata
);

  axi_writer #(
            .C_M_AXI_ADDR_WIDTH  ( C_M_AXI_ADDR_WIDTH ) ,
            .C_M_AXI_DATA_WIDTH  ( C_M_AXI_DATA_WIDTH ) ,
            .C_XFER_SIZE_WIDTH   ( C_XFER_SIZE_WIDTH  ) ,
            .C_MAX_OUTSTANDING   ( C_MAX_OUTSTANDING  ) ,
            .C_INCLUDE_DATA_FIFO ( C_INCLUDE_DATA_FIFO)
          )
          inst_axi_writer (
            .aclk                    ( aclk                   ) ,
            .areset                  ( areset                 ) ,
            .ctrl_start              ( ctrl_start             ) ,
            .ctrl_done               ( ctrl_done              ) ,
            .ctrl_addr_offset        ( ctrl_addr_offset       ) ,
            .ctrl_xfer_size_in_bytes ( ctrl_xfer_size_in_bytes) ,
            .m_axi_awvalid           ( m_axi_awvalid) ,
            .m_axi_awready           ( m_axi_awready) ,
            .m_axi_awaddr            ( m_axi_awaddr ) ,
            .m_axi_awlen             ( m_axi_awlen  ) ,
            .m_axi_wvalid            ( m_axi_wvalid ) ,
            .m_axi_wready            ( m_axi_wready ) ,
            .m_axi_wdata             ( m_axi_wdata  ) ,
            .m_axi_wstrb             ( m_axi_wstrb  ) ,
            .m_axi_wlast             ( m_axi_wlast  ) ,
            .m_axi_bvalid            ( m_axi_bvalid ) ,
            .m_axi_bready            ( m_axi_bready ) ,
            .s_axis_aclk             ( s_axis_aclk  ) ,
            .s_axis_areset           ( s_axis_areset) ,
            .s_axis_tvalid           (s_axis_tvalid ) ,
            .s_axis_tready           (s_axis_tready ) ,
            .s_axis_tdata            (s_axis_tdata  )
          );

endmodule



module m_accelerator
(
  input clk,
  input rst,
  input start,
  input [32-1:0] acc_user_done_rd_data,
  input [32-1:0] acc_user_done_wr_data,
  output [32-1:0] acc_user_request_read,
  input [32-1:0] acc_user_read_data_valid,
  input [8192-1:0] acc_user_read_data,
  input [32-1:0] acc_user_available_write,
  output [32-1:0] acc_user_request_write,
  output [8192-1:0] acc_user_write_data,
  output acc_user_done
);
  
  reg [32-1:0] request_read;
  reg [32-1:0] request_write;
  reg [8192-1:0] write_data;
  reg [32-1:0] done_rd_data;
  reg [32-1:0] done_wr_data;
  reg done;
  
  assign acc_user_done = done;
  assign acc_user_request_read = request_read;
  assign acc_user_request_write = request_write;
  assign acc_user_write_data = write_data;
  
  always @(posedge clk)begin
      if(rst)begin
          done <= 0;
          done_rd_data <= 0;
          done_wr_data <= 0;
      end
      else begin
        done_rd_data <= acc_user_done_rd_data;
        done_wr_data <= acc_user_done_wr_data;
        done <= &{done_rd_data,done_wr_data};
      end
  end
  
  integer i;
 
    always @(posedge clk)begin
        if(rst)begin
          request_write <= 0;
          request_read <= 0;
        end
        else begin
          write_data <= acc_user_read_data;
          request_write <= 0;
          request_read <= 0;
          for(i=0;i < 32;i =  i + 1)begin
            if(acc_user_available_write[i] & acc_user_read_data_valid[i])begin
               request_write[i] <= 1;
               request_read[i] <= 1;
            end
          end
        end
    end
    
    reg [32-1:0]count_rd[0:32-1];
    reg [32-1:0]count_wr[0:32-1];
  
    always @(posedge clk)begin
      if(rst)begin
         for(i=0;i < 32;i =  i + 1)begin
           count_rd[i] <= 0;
           count_wr[i] <= 0;
        end
      end else begin
       for(i=0;i < 32;i =  i + 1)begin
           if(request_read[i])begin
             count_rd[i] <= count_rd[i]+1;
           end
           if(request_write[i])begin
             count_wr[i] <= count_wr[i]+1;
           end
       end 
      end
    end
  
endmodule
